/* Description : This verilog file tends to build the FFT Block using the following blocks : */
/* RAM , MUX , Butterfly Column , Registers and Controller  */
/* Authors : Basma Walid and Mohammed Abd el Nasser - Preprocessing Team */

/* NOTE : Number of Registers used is 256 . However , Every two registers are connected to the same enable */

module FFT_Time_Share_Top_Module #(
	parameter BITS = 16 ,						/* Number of bits of the data(inputs and outputs) */
	parameter SEL_BITS = 7 ,					/* Number of bits of the MUX Selection lines */
	parameter ADDRESS_BITS = 2 ,				/* Number of bits of the memory address bus */
	parameter NUMBER_OF_LOCATIONS = 4 ,			/* Number of locations of the memory*/
	parameter NUMBER_OF_ENABLE_BITS = 128,		/* Number of enable bits of the Registers used */
	parameter NUMBER_OF_MEM = 32 				/* Number of Memory instances i.e Memory Enables */
)
(
	input wire ready_inputs ,
	input wire clk ,
	input wire rst ,
	input wire [BITS-1:0] x0_r ,
	input wire [BITS-1:0] x0_i ,
	input wire [BITS-1:0] x1_r ,
    input wire [BITS-1:0] x1_i ,
    input wire [BITS-1:0] x2_r ,
    input wire [BITS-1:0] x2_i ,
    input wire [BITS-1:0] x3_r ,
    input wire [BITS-1:0] x3_i ,
    input wire [BITS-1:0] x4_r ,
    input wire [BITS-1:0] x4_i ,
    input wire [BITS-1:0] x5_r ,
    input wire [BITS-1:0] x5_i ,
    input wire [BITS-1:0] x6_r ,
    input wire [BITS-1:0] x6_i ,
    input wire [BITS-1:0] x7_r ,
    input wire [BITS-1:0] x7_i ,
    input wire [BITS-1:0] x8_r ,
    input wire [BITS-1:0] x8_i ,
    input wire [BITS-1:0] x9_r ,
    input wire [BITS-1:0] x9_i ,
    input wire [BITS-1:0] x10_r ,
    input wire [BITS-1:0] x10_i ,
    input wire [BITS-1:0] x11_r ,
    input wire [BITS-1:0] x11_i ,
    input wire [BITS-1:0] x12_r ,
    input wire [BITS-1:0] x12_i ,
    input wire [BITS-1:0] x13_r ,
    input wire [BITS-1:0] x13_i ,
    input wire [BITS-1:0] x14_r ,
    input wire [BITS-1:0] x14_i ,
    input wire [BITS-1:0] x15_r ,
    input wire [BITS-1:0] x15_i ,
    input wire [BITS-1:0] x16_r ,
    input wire [BITS-1:0] x16_i ,
    input wire [BITS-1:0] x17_r ,
    input wire [BITS-1:0] x17_i ,
    input wire [BITS-1:0] x18_r ,
    input wire [BITS-1:0] x18_i ,
    input wire [BITS-1:0] x19_r ,
    input wire [BITS-1:0] x19_i ,
    input wire [BITS-1:0] x20_r ,
    input wire [BITS-1:0] x20_i ,
    input wire [BITS-1:0] x21_r ,
    input wire [BITS-1:0] x21_i ,
    input wire [BITS-1:0] x22_r ,
    input wire [BITS-1:0] x22_i ,
    input wire [BITS-1:0] x23_r ,
    input wire [BITS-1:0] x23_i ,
    input wire [BITS-1:0] x24_r ,
    input wire [BITS-1:0] x24_i ,
    input wire [BITS-1:0] x25_r ,
    input wire [BITS-1:0] x25_i ,
    input wire [BITS-1:0] x26_r ,
    input wire [BITS-1:0] x26_i ,
    input wire [BITS-1:0] x27_r ,
    input wire [BITS-1:0] x27_i ,
    input wire [BITS-1:0] x28_r ,
    input wire [BITS-1:0] x28_i ,
    input wire [BITS-1:0] x29_r ,
    input wire [BITS-1:0] x29_i ,
    input wire [BITS-1:0] x30_r ,
    input wire [BITS-1:0] x30_i ,
    input wire [BITS-1:0] x31_r ,
    input wire [BITS-1:0] x31_i ,
    input wire [BITS-1:0] x32_r ,
    input wire [BITS-1:0] x32_i ,
    input wire [BITS-1:0] x33_r ,
    input wire [BITS-1:0] x33_i ,
    input wire [BITS-1:0] x34_r ,
    input wire [BITS-1:0] x34_i ,
    input wire [BITS-1:0] x35_r ,
    input wire [BITS-1:0] x35_i ,
    input wire [BITS-1:0] x36_r ,
    input wire [BITS-1:0] x36_i ,
    input wire [BITS-1:0] x37_r ,
    input wire [BITS-1:0] x37_i ,
    input wire [BITS-1:0] x38_r ,
    input wire [BITS-1:0] x38_i ,
    input wire [BITS-1:0] x39_r ,
    input wire [BITS-1:0] x39_i ,
    input wire [BITS-1:0] x40_r ,
    input wire [BITS-1:0] x40_i ,
    input wire [BITS-1:0] x41_r ,
    input wire [BITS-1:0] x41_i ,
    input wire [BITS-1:0] x42_r ,
    input wire [BITS-1:0] x42_i ,
    input wire [BITS-1:0] x43_r ,
    input wire [BITS-1:0] x43_i ,
    input wire [BITS-1:0] x44_r ,
    input wire [BITS-1:0] x44_i ,
    input wire [BITS-1:0] x45_r ,
    input wire [BITS-1:0] x45_i ,
    input wire [BITS-1:0] x46_r ,
    input wire [BITS-1:0] x46_i ,
    input wire [BITS-1:0] x47_r ,
    input wire [BITS-1:0] x47_i ,
    input wire [BITS-1:0] x48_r ,
    input wire [BITS-1:0] x48_i ,
    input wire [BITS-1:0] x49_r ,
    input wire [BITS-1:0] x49_i ,
    input wire [BITS-1:0] x50_r ,
    input wire [BITS-1:0] x50_i ,
    input wire [BITS-1:0] x51_r ,
    input wire [BITS-1:0] x51_i ,
    input wire [BITS-1:0] x52_r ,
    input wire [BITS-1:0] x52_i ,
    input wire [BITS-1:0] x53_r ,
    input wire [BITS-1:0] x53_i ,
    input wire [BITS-1:0] x54_r ,
    input wire [BITS-1:0] x54_i ,
    input wire [BITS-1:0] x55_r ,
    input wire [BITS-1:0] x55_i ,
    input wire [BITS-1:0] x56_r ,
    input wire [BITS-1:0] x56_i ,
    input wire [BITS-1:0] x57_r ,
    input wire [BITS-1:0] x57_i ,
    input wire [BITS-1:0] x58_r ,
    input wire [BITS-1:0] x58_i ,
    input wire [BITS-1:0] x59_r ,
    input wire [BITS-1:0] x59_i ,
    input wire [BITS-1:0] x60_r ,
    input wire [BITS-1:0] x60_i ,
    input wire [BITS-1:0] x61_r ,
    input wire [BITS-1:0] x61_i ,
    input wire [BITS-1:0] x62_r ,
    input wire [BITS-1:0] x62_i ,
    input wire [BITS-1:0] x63_r ,
    input wire [BITS-1:0] x63_i ,
    input wire [BITS-1:0] x64_r ,
    input wire [BITS-1:0] x64_i ,
    input wire [BITS-1:0] x65_r ,
    input wire [BITS-1:0] x65_i ,
    input wire [BITS-1:0] x66_r ,
    input wire [BITS-1:0] x66_i ,
    input wire [BITS-1:0] x67_r ,
    input wire [BITS-1:0] x67_i ,
    input wire [BITS-1:0] x68_r ,
    input wire [BITS-1:0] x68_i ,
    input wire [BITS-1:0] x69_r ,
    input wire [BITS-1:0] x69_i ,
    input wire [BITS-1:0] x70_r ,
    input wire [BITS-1:0] x70_i ,
    input wire [BITS-1:0] x71_r ,
    input wire [BITS-1:0] x71_i ,
    input wire [BITS-1:0] x72_r ,
    input wire [BITS-1:0] x72_i ,
    input wire [BITS-1:0] x73_r ,
    input wire [BITS-1:0] x73_i ,
    input wire [BITS-1:0] x74_r ,
    input wire [BITS-1:0] x74_i ,
    input wire [BITS-1:0] x75_r ,
    input wire [BITS-1:0] x75_i ,
    input wire [BITS-1:0] x76_r ,
    input wire [BITS-1:0] x76_i ,
    input wire [BITS-1:0] x77_r ,
    input wire [BITS-1:0] x77_i ,
    input wire [BITS-1:0] x78_r ,
    input wire [BITS-1:0] x78_i ,
    input wire [BITS-1:0] x79_r ,
    input wire [BITS-1:0] x79_i ,
    input wire [BITS-1:0] x80_r ,
    input wire [BITS-1:0] x80_i ,
    input wire [BITS-1:0] x81_r ,
    input wire [BITS-1:0] x81_i ,
    input wire [BITS-1:0] x82_r ,
    input wire [BITS-1:0] x82_i ,
    input wire [BITS-1:0] x83_r ,
    input wire [BITS-1:0] x83_i ,
    input wire [BITS-1:0] x84_r ,
    input wire [BITS-1:0] x84_i ,
    input wire [BITS-1:0] x85_r ,
    input wire [BITS-1:0] x85_i ,
    input wire [BITS-1:0] x86_r ,
    input wire [BITS-1:0] x86_i ,
    input wire [BITS-1:0] x87_r ,
    input wire [BITS-1:0] x87_i ,
    input wire [BITS-1:0] x88_r ,
    input wire [BITS-1:0] x88_i ,
    input wire [BITS-1:0] x89_r ,
    input wire [BITS-1:0] x89_i ,
    input wire [BITS-1:0] x90_r ,
    input wire [BITS-1:0] x90_i ,
    input wire [BITS-1:0] x91_r ,
    input wire [BITS-1:0] x91_i ,
    input wire [BITS-1:0] x92_r ,
    input wire [BITS-1:0] x92_i ,
    input wire [BITS-1:0] x93_r ,
    input wire [BITS-1:0] x93_i ,
    input wire [BITS-1:0] x94_r ,
    input wire [BITS-1:0] x94_i ,
    input wire [BITS-1:0] x95_r ,
    input wire [BITS-1:0] x95_i ,
    input wire [BITS-1:0] x96_r ,
    input wire [BITS-1:0] x96_i ,
    input wire [BITS-1:0] x97_r ,
    input wire [BITS-1:0] x97_i ,
    input wire [BITS-1:0] x98_r ,
    input wire [BITS-1:0] x98_i ,
    input wire [BITS-1:0] x99_r ,
    input wire [BITS-1:0] x99_i ,
    input wire [BITS-1:0] x100_r ,
    input wire [BITS-1:0] x100_i ,
    input wire [BITS-1:0] x101_r ,
    input wire [BITS-1:0] x101_i ,
    input wire [BITS-1:0] x102_r ,
    input wire [BITS-1:0] x102_i ,
    input wire [BITS-1:0] x103_r ,
    input wire [BITS-1:0] x103_i ,
    input wire [BITS-1:0] x104_r ,
    input wire [BITS-1:0] x104_i ,
    input wire [BITS-1:0] x105_r ,
    input wire [BITS-1:0] x105_i ,
    input wire [BITS-1:0] x106_r ,
    input wire [BITS-1:0] x106_i ,
    input wire [BITS-1:0] x107_r ,
    input wire [BITS-1:0] x107_i ,
    input wire [BITS-1:0] x108_r ,
    input wire [BITS-1:0] x108_i ,
    input wire [BITS-1:0] x109_r ,
    input wire [BITS-1:0] x109_i ,
    input wire [BITS-1:0] x110_r ,
    input wire [BITS-1:0] x110_i ,
    input wire [BITS-1:0] x111_r ,
    input wire [BITS-1:0] x111_i ,
    input wire [BITS-1:0] x112_r ,
    input wire [BITS-1:0] x112_i ,
    input wire [BITS-1:0] x113_r ,
    input wire [BITS-1:0] x113_i ,
    input wire [BITS-1:0] x114_r ,
    input wire [BITS-1:0] x114_i ,
    input wire [BITS-1:0] x115_r ,
    input wire [BITS-1:0] x115_i ,
    input wire [BITS-1:0] x116_r ,
    input wire [BITS-1:0] x116_i ,
    input wire [BITS-1:0] x117_r ,
    input wire [BITS-1:0] x117_i ,
    input wire [BITS-1:0] x118_r ,
    input wire [BITS-1:0] x118_i ,
    input wire [BITS-1:0] x119_r ,
    input wire [BITS-1:0] x119_i ,
    input wire [BITS-1:0] x120_r ,
    input wire [BITS-1:0] x120_i ,
    input wire [BITS-1:0] x121_r ,
    input wire [BITS-1:0] x121_i ,
    input wire [BITS-1:0] x122_r ,
    input wire [BITS-1:0] x122_i ,
    input wire [BITS-1:0] x123_r ,
    input wire [BITS-1:0] x123_i ,
    input wire [BITS-1:0] x124_r ,
    input wire [BITS-1:0] x124_i ,
    input wire [BITS-1:0] x125_r ,
    input wire [BITS-1:0] x125_i ,
    input wire [BITS-1:0] x126_r ,
    input wire [BITS-1:0] x126_i ,
    input wire [BITS-1:0] x127_r ,
    input wire [BITS-1:0] x127_i ,
	
	output wire correct ,
	output wire [BITS-1:0] X0_r ,
    output wire [BITS-1:0] X0_i ,
    output wire [BITS-1:0] X1_r ,
    output wire [BITS-1:0] X1_i ,
    output wire [BITS-1:0] X2_r ,
    output wire [BITS-1:0] X2_i ,
    output wire [BITS-1:0] X3_r ,
    output wire [BITS-1:0] X3_i ,
    output wire [BITS-1:0] X4_r ,
    output wire [BITS-1:0] X4_i ,
    output wire [BITS-1:0] X5_r ,
    output wire [BITS-1:0] X5_i ,
    output wire [BITS-1:0] X6_r ,
    output wire [BITS-1:0] X6_i ,
    output wire [BITS-1:0] X7_r ,
    output wire [BITS-1:0] X7_i ,
    output wire [BITS-1:0] X8_r ,
    output wire [BITS-1:0] X8_i ,
    output wire [BITS-1:0] X9_r ,
    output wire [BITS-1:0] X9_i ,
    output wire [BITS-1:0] X10_r ,
    output wire [BITS-1:0] X10_i ,
    output wire [BITS-1:0] X11_r ,
    output wire [BITS-1:0] X11_i ,
    output wire [BITS-1:0] X12_r ,
    output wire [BITS-1:0] X12_i ,
    output wire [BITS-1:0] X13_r ,
    output wire [BITS-1:0] X13_i ,
    output wire [BITS-1:0] X14_r ,
    output wire [BITS-1:0] X14_i ,
    output wire [BITS-1:0] X15_r ,
    output wire [BITS-1:0] X15_i ,
    output wire [BITS-1:0] X16_r ,
    output wire [BITS-1:0] X16_i ,
    output wire [BITS-1:0] X17_r ,
    output wire [BITS-1:0] X17_i ,
    output wire [BITS-1:0] X18_r ,
    output wire [BITS-1:0] X18_i ,
    output wire [BITS-1:0] X19_r ,
    output wire [BITS-1:0] X19_i ,
    output wire [BITS-1:0] X20_r ,
    output wire [BITS-1:0] X20_i ,
    output wire [BITS-1:0] X21_r ,
    output wire [BITS-1:0] X21_i ,
    output wire [BITS-1:0] X22_r ,
    output wire [BITS-1:0] X22_i ,
    output wire [BITS-1:0] X23_r ,
    output wire [BITS-1:0] X23_i ,
    output wire [BITS-1:0] X24_r ,
    output wire [BITS-1:0] X24_i ,
    output wire [BITS-1:0] X25_r ,
    output wire [BITS-1:0] X25_i ,
    output wire [BITS-1:0] X26_r ,
    output wire [BITS-1:0] X26_i ,
    output wire [BITS-1:0] X27_r ,
    output wire [BITS-1:0] X27_i ,
    output wire [BITS-1:0] X28_r ,
    output wire [BITS-1:0] X28_i ,
    output wire [BITS-1:0] X29_r ,
    output wire [BITS-1:0] X29_i ,
    output wire [BITS-1:0] X30_r ,
    output wire [BITS-1:0] X30_i ,
    output wire [BITS-1:0] X31_r ,
    output wire [BITS-1:0] X31_i ,
    output wire [BITS-1:0] X32_r ,
    output wire [BITS-1:0] X32_i ,
    output wire [BITS-1:0] X33_r ,
    output wire [BITS-1:0] X33_i ,
    output wire [BITS-1:0] X34_r ,
    output wire [BITS-1:0] X34_i ,
    output wire [BITS-1:0] X35_r ,
    output wire [BITS-1:0] X35_i ,
    output wire [BITS-1:0] X36_r ,
    output wire [BITS-1:0] X36_i ,
    output wire [BITS-1:0] X37_r ,
    output wire [BITS-1:0] X37_i ,
    output wire [BITS-1:0] X38_r ,
    output wire [BITS-1:0] X38_i ,
    output wire [BITS-1:0] X39_r ,
    output wire [BITS-1:0] X39_i ,
    output wire [BITS-1:0] X40_r ,
    output wire [BITS-1:0] X40_i ,
    output wire [BITS-1:0] X41_r ,
    output wire [BITS-1:0] X41_i ,
    output wire [BITS-1:0] X42_r ,
    output wire [BITS-1:0] X42_i ,
    output wire [BITS-1:0] X43_r ,
    output wire [BITS-1:0] X43_i ,
    output wire [BITS-1:0] X44_r ,
    output wire [BITS-1:0] X44_i ,
    output wire [BITS-1:0] X45_r ,
    output wire [BITS-1:0] X45_i ,
    output wire [BITS-1:0] X46_r ,
    output wire [BITS-1:0] X46_i ,
    output wire [BITS-1:0] X47_r ,
    output wire [BITS-1:0] X47_i ,
    output wire [BITS-1:0] X48_r ,
    output wire [BITS-1:0] X48_i ,
    output wire [BITS-1:0] X49_r ,
    output wire [BITS-1:0] X49_i ,
    output wire [BITS-1:0] X50_r ,
    output wire [BITS-1:0] X50_i ,
    output wire [BITS-1:0] X51_r ,
    output wire [BITS-1:0] X51_i ,
    output wire [BITS-1:0] X52_r ,
    output wire [BITS-1:0] X52_i ,
    output wire [BITS-1:0] X53_r ,
    output wire [BITS-1:0] X53_i ,
    output wire [BITS-1:0] X54_r ,
    output wire [BITS-1:0] X54_i ,
    output wire [BITS-1:0] X55_r ,
    output wire [BITS-1:0] X55_i ,
    output wire [BITS-1:0] X56_r ,
    output wire [BITS-1:0] X56_i ,
    output wire [BITS-1:0] X57_r ,
    output wire [BITS-1:0] X57_i ,
    output wire [BITS-1:0] X58_r ,
    output wire [BITS-1:0] X58_i ,
    output wire [BITS-1:0] X59_r ,
    output wire [BITS-1:0] X59_i ,
    output wire [BITS-1:0] X60_r ,
    output wire [BITS-1:0] X60_i ,
    output wire [BITS-1:0] X61_r ,
    output wire [BITS-1:0] X61_i ,
    output wire [BITS-1:0] X62_r ,
    output wire [BITS-1:0] X62_i ,
    output wire [BITS-1:0] X63_r ,
    output wire [BITS-1:0] X63_i ,
    output wire [BITS-1:0] X64_r ,
    output wire [BITS-1:0] X64_i ,
    output wire [BITS-1:0] X65_r ,
    output wire [BITS-1:0] X65_i ,
    output wire [BITS-1:0] X66_r ,
    output wire [BITS-1:0] X66_i ,
    output wire [BITS-1:0] X67_r ,
    output wire [BITS-1:0] X67_i ,
    output wire [BITS-1:0] X68_r ,
    output wire [BITS-1:0] X68_i ,
    output wire [BITS-1:0] X69_r ,
    output wire [BITS-1:0] X69_i ,
    output wire [BITS-1:0] X70_r ,
    output wire [BITS-1:0] X70_i ,
    output wire [BITS-1:0] X71_r ,
    output wire [BITS-1:0] X71_i ,
    output wire [BITS-1:0] X72_r ,
    output wire [BITS-1:0] X72_i ,
    output wire [BITS-1:0] X73_r ,
    output wire [BITS-1:0] X73_i ,
    output wire [BITS-1:0] X74_r ,
    output wire [BITS-1:0] X74_i ,
    output wire [BITS-1:0] X75_r ,
    output wire [BITS-1:0] X75_i ,
    output wire [BITS-1:0] X76_r ,
    output wire [BITS-1:0] X76_i ,
    output wire [BITS-1:0] X77_r ,
    output wire [BITS-1:0] X77_i ,
    output wire [BITS-1:0] X78_r ,
    output wire [BITS-1:0] X78_i ,
    output wire [BITS-1:0] X79_r ,
    output wire [BITS-1:0] X79_i ,
    output wire [BITS-1:0] X80_r ,
    output wire [BITS-1:0] X80_i ,
    output wire [BITS-1:0] X81_r ,
    output wire [BITS-1:0] X81_i ,
    output wire [BITS-1:0] X82_r ,
    output wire [BITS-1:0] X82_i ,
    output wire [BITS-1:0] X83_r ,
    output wire [BITS-1:0] X83_i ,
    output wire [BITS-1:0] X84_r ,
    output wire [BITS-1:0] X84_i ,
    output wire [BITS-1:0] X85_r ,
    output wire [BITS-1:0] X85_i ,
    output wire [BITS-1:0] X86_r ,
    output wire [BITS-1:0] X86_i ,
    output wire [BITS-1:0] X87_r ,
    output wire [BITS-1:0] X87_i ,
    output wire [BITS-1:0] X88_r ,
    output wire [BITS-1:0] X88_i ,
    output wire [BITS-1:0] X89_r ,
    output wire [BITS-1:0] X89_i ,
    output wire [BITS-1:0] X90_r ,
    output wire [BITS-1:0] X90_i ,
    output wire [BITS-1:0] X91_r ,
    output wire [BITS-1:0] X91_i ,
    output wire [BITS-1:0] X92_r ,
    output wire [BITS-1:0] X92_i ,
    output wire [BITS-1:0] X93_r ,
    output wire [BITS-1:0] X93_i ,
    output wire [BITS-1:0] X94_r ,
    output wire [BITS-1:0] X94_i ,
    output wire [BITS-1:0] X95_r ,
    output wire [BITS-1:0] X95_i ,
    output wire [BITS-1:0] X96_r ,
    output wire [BITS-1:0] X96_i ,
    output wire [BITS-1:0] X97_r ,
    output wire [BITS-1:0] X97_i ,
    output wire [BITS-1:0] X98_r ,
    output wire [BITS-1:0] X98_i ,
    output wire [BITS-1:0] X99_r ,
    output wire [BITS-1:0] X99_i ,
    output wire [BITS-1:0] X100_r ,
    output wire [BITS-1:0] X100_i ,
    output wire [BITS-1:0] X101_r ,
    output wire [BITS-1:0] X101_i ,
    output wire [BITS-1:0] X102_r ,
    output wire [BITS-1:0] X102_i ,
    output wire [BITS-1:0] X103_r ,
    output wire [BITS-1:0] X103_i ,
    output wire [BITS-1:0] X104_r ,
    output wire [BITS-1:0] X104_i ,
    output wire [BITS-1:0] X105_r ,
    output wire [BITS-1:0] X105_i ,
    output wire [BITS-1:0] X106_r ,
    output wire [BITS-1:0] X106_i ,
    output wire [BITS-1:0] X107_r ,
    output wire [BITS-1:0] X107_i ,
    output wire [BITS-1:0] X108_r ,
    output wire [BITS-1:0] X108_i ,
    output wire [BITS-1:0] X109_r ,
    output wire [BITS-1:0] X109_i ,
    output wire [BITS-1:0] X110_r ,
    output wire [BITS-1:0] X110_i ,
    output wire [BITS-1:0] X111_r ,
    output wire [BITS-1:0] X111_i ,
    output wire [BITS-1:0] X112_r ,
    output wire [BITS-1:0] X112_i ,
    output wire [BITS-1:0] X113_r ,
    output wire [BITS-1:0] X113_i ,
    output wire [BITS-1:0] X114_r ,
    output wire [BITS-1:0] X114_i ,
    output wire [BITS-1:0] X115_r ,
    output wire [BITS-1:0] X115_i ,
    output wire [BITS-1:0] X116_r ,
    output wire [BITS-1:0] X116_i ,
    output wire [BITS-1:0] X117_r ,
    output wire [BITS-1:0] X117_i ,
    output wire [BITS-1:0] X118_r ,
    output wire [BITS-1:0] X118_i ,
    output wire [BITS-1:0] X119_r ,
    output wire [BITS-1:0] X119_i ,
    output wire [BITS-1:0] X120_r ,
    output wire [BITS-1:0] X120_i ,
    output wire [BITS-1:0] X121_r ,
    output wire [BITS-1:0] X121_i ,
    output wire [BITS-1:0] X122_r ,
    output wire [BITS-1:0] X122_i ,
    output wire [BITS-1:0] X123_r ,
    output wire [BITS-1:0] X123_i ,
    output wire [BITS-1:0] X124_r ,
    output wire [BITS-1:0] X124_i ,
    output wire [BITS-1:0] X125_r ,
    output wire [BITS-1:0] X125_i ,
    output wire [BITS-1:0] X126_r ,
    output wire [BITS-1:0] X126_i ,
    output wire [BITS-1:0] X127_r ,
    output wire [BITS-1:0] X127_i 
);

/* Internal Signals */

/* CONTROLLER */
/* Outputs */
wire [SEL_BITS-1:0]  sel_output_mux_0 ; /*Input to MUX_0. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_1 ; /*Input to MUX_1. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_2 ; /*Input to MUX_2. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_3 ; /*Input to MUX_3. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_4 ; /*Input to MUX_4. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_5 ; /*Input to MUX_5. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_6 ; /*Input to MUX_6. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_7 ; /*Input to MUX_7. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_8 ; /*Input to MUX_8. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_9 ; /*Input to MUX_9. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_10 ; /*Input to MUX_10. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_11 ; /*Input to MUX_11. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_12 ; /*Input to MUX_12. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_13 ; /*Input to MUX_13. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_14 ; /*Input to MUX_14. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_15 ; /*Input to MUX_15. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_16 ; /*Input to MUX_16. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_17 ; /*Input to MUX_17. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_18 ; /*Input to MUX_18. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_19 ; /*Input to MUX_19. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_20 ; /*Input to MUX_20. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_21 ; /*Input to MUX_21. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_22 ; /*Input to MUX_22. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_23 ; /*Input to MUX_23. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_24 ; /*Input to MUX_24. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_25 ; /*Input to MUX_25. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_26 ; /*Input to MUX_26. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_27 ; /*Input to MUX_27. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_28 ; /*Input to MUX_28. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_29 ; /*Input to MUX_29. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_30 ; /*Input to MUX_30. Output of Controller */
wire [SEL_BITS-1:0]  sel_output_mux_31 ; /*Input to MUX_31. Output of Controller */

wire [NUMBER_OF_ENABLE_BITS-1:0] reg_en; /*Input to the Registers. Output of Controller */
wire [63:0] twiddle_reg_en;              /*Input to the twiddle Registers. Output of Controller */
wire [4:0] ROM_addr ;                    /*Input to the twiddle ROM. Output of Controller */
wire [ADDRESS_BITS-1:0] read_address ;   /*Input to the Memory. Output of Controller */
wire [ADDRESS_BITS-1:0] write_address ;	 /*Input to the Memory. Output of Controller */
wire [NUMBER_OF_MEM-1:0] mem_write_enable ; /*Input to the Memory. Output of Controller */
wire [1:0]  sel_output_4x1 ;

/* Butterfly Column Internal Signals */
/* Inputs */

/* Outputs */
wire [BITS-1:0] s0_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s0_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s1_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s1_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s2_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s2_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s3_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s3_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s4_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s4_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s5_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s5_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s6_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s6_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s7_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s7_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s8_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s8_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s9_r ; 					/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s9_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s10_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s10_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s11_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s11_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s12_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s12_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s13_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s13_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s14_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s14_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s15_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s15_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s16_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s16_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s17_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s17_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s18_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s18_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s19_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s19_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s20_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s20_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s21_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s21_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s22_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s22_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s23_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s23_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s24_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s24_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s25_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s25_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s26_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s26_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s27_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s27_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s28_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s28_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s29_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s29_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s30_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s30_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s31_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s31_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s32_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s32_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s33_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s33_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s34_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s34_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s35_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s35_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s36_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s36_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s37_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s37_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s38_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s38_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s39_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s39_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s40_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s40_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s41_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s41_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s42_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s42_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s43_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s43_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s44_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s44_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s45_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s45_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s46_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s46_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s47_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s47_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s48_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s48_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s49_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s49_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s50_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s50_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s51_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s51_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s52_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s52_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s53_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s53_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s54_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s54_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s55_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s55_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s56_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s56_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s57_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s57_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s58_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s58_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s59_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s59_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s60_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s60_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s61_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s61_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s62_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s62_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s63_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s63_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s64_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s64_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s65_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s65_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s66_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s66_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s67_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s67_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s68_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s68_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s69_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s69_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s70_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s70_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s71_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s71_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s72_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s72_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s73_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s73_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s74_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s74_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s75_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s75_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s76_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s76_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s77_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s77_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s78_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s78_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s79_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s79_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s80_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s80_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s81_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s81_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s82_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s82_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s83_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s83_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s84_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s84_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s85_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s85_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s86_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s86_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s87_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s87_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s88_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s88_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s89_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s89_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s90_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s90_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s91_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s91_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s92_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s92_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s93_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s93_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s94_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s94_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s95_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s95_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s96_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s96_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s97_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s97_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s98_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s98_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s99_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s99_i ;					/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s100_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s100_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s101_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s101_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s102_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s102_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s103_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s103_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s104_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s104_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s105_r ;				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s105_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s106_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s106_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s107_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s107_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s108_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s108_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s109_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s109_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s110_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s110_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s111_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s111_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s112_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s112_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s113_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s113_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s114_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s114_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s115_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s115_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s116_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s116_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s117_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s117_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s118_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s118_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s119_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s119_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s120_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s120_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s121_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s121_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s122_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s122_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s123_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s123_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s124_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s124_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s125_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s125_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s126_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s126_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s127_r ; 				/* Input to all instances of MUX_REAL_MEMORY. Output of Butterfly Column */ 
wire [BITS-1:0] s127_i ;				/* Input to all instances of MUX_IMG_MEMORY. Output of Butterfly Column */


/* REAL MEMORY */
/* Inputs */
wire [BITS-1:0] mux_2_1_0_output_real ;    /* Input to Memory . Output of 2x1 U0_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_1_output_real ;    /* Input to Memory . Output of 2x1 U1_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_2_output_real ;    /* Input to Memory . Output of 2x1 U2_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_3_output_real ;    /* Input to Memory . Output of 2x1 U3_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_4_output_real ;    /* Input to Memory . Output of 2x1 U4_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_5_output_real ;    /* Input to Memory . Output of 2x1 U5_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_6_output_real ;    /* Input to Memory . Output of 2x1 U6_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_7_output_real ;    /* Input to Memory . Output of 2x1 U7_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_8_output_real ;    /* Input to Memory . Output of 2x1 U8_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_9_output_real ;    /* Input to Memory . Output of 2x1 U9_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_10_output_real ;    /* Input to Memory . Output of 2x1 U10_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_11_output_real ;    /* Input to Memory . Output of 2x1 U11_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_12_output_real ;    /* Input to Memory . Output of 2x1 U12_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_13_output_real ;    /* Input to Memory . Output of 2x1 U13_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_14_output_real ;    /* Input to Memory . Output of 2x1 U14_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_15_output_real ;    /* Input to Memory . Output of 2x1 U15_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_16_output_real ;    /* Input to Memory . Output of 2x1 U16_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_17_output_real ;    /* Input to Memory . Output of 2x1 U17_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_18_output_real ;    /* Input to Memory . Output of 2x1 U18_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_19_output_real ;    /* Input to Memory . Output of 2x1 U19_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_20_output_real ;    /* Input to Memory . Output of 2x1 U20_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_21_output_real ;    /* Input to Memory . Output of 2x1 U21_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_22_output_real ;    /* Input to Memory . Output of 2x1 U22_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_23_output_real ;    /* Input to Memory . Output of 2x1 U23_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_24_output_real ;    /* Input to Memory . Output of 2x1 U24_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_25_output_real ;    /* Input to Memory . Output of 2x1 U25_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_26_output_real ;    /* Input to Memory . Output of 2x1 U26_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_27_output_real ;    /* Input to Memory . Output of 2x1 U27_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_28_output_real ;    /* Input to Memory . Output of 2x1 U28_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_29_output_real ;    /* Input to Memory . Output of 2x1 U29_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_30_output_real ;    /* Input to Memory . Output of 2x1 U30_REAL_MUX_2_1 */
wire [BITS-1:0] mux_2_1_31_output_real ;    /* Input to Memory . Output of 2x1 U31_REAL_MUX_2_1 */


/* Outputs */
wire [BITS-1:0] memory_real_output_0 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_1 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_2 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_3 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_4 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_5 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_6 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_7 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_8 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_9 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_10 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_11 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_12 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_13 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_14 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_15 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_16 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_17 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_18 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_19 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_20 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_21 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_22 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_23 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_24 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_25 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_26 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_27 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_28 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_29 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_30 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_real_output_31 ;  /* Output of Memory . Input to Registers */

/* MUX 2x1 */
wire [BITS-1:0] mux_0_output_real ;		/* Input to 2x1 U0_REAL_MUX_2_1 . Output of 128x1 U0_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_1_output_real ;		/* Input to 2x1 U1_REAL_MUX_2_1 . Output of 128x1 U1_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_2_output_real ;		/* Input to 2x1 U2_REAL_MUX_2_1 . Output of 128x1 U2_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_3_output_real ;		/* Input to 2x1 U3_REAL_MUX_2_1 . Output of 128x1 U3_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_4_output_real ;		/* Input to 2x1 U4_REAL_MUX_2_1 . Output of 128x1 U4_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_5_output_real ;		/* Input to 2x1 U5_REAL_MUX_2_1 . Output of 128x1 U5_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_6_output_real ;		/* Input to 2x1 U6_REAL_MUX_2_1 . Output of 128x1 U6_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_7_output_real ;		/* Input to 2x1 U7_REAL_MUX_2_1 . Output of 128x1 U7_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_8_output_real ;		/* Input to 2x1 U8_REAL_MUX_2_1 . Output of 128x1 U8_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_9_output_real ;		/* Input to 2x1 U9_REAL_MUX_2_1 . Output of 128x1 U9_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_10_output_real ;	/* Input to 2x1 U10_REAL_MUX_2_1 . Output of 128x1 U10_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_11_output_real ;	/* Input to 2x1 U11_REAL_MUX_2_1 . Output of 128x1 U11_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_12_output_real ;	/* Input to 2x1 U12_REAL_MUX_2_1 . Output of 128x1 U12_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_13_output_real ;	/* Input to 2x1 U13_REAL_MUX_2_1 . Output of 128x1 U13_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_14_output_real ;	/* Input to 2x1 U14_REAL_MUX_2_1 . Output of 128x1 U14_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_15_output_real ;	/* Input to 2x1 U15_REAL_MUX_2_1 . Output of 128x1 U15_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_16_output_real ;	/* Input to 2x1 U16_REAL_MUX_2_1 . Output of 128x1 U16_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_17_output_real ;	/* Input to 2x1 U17_REAL_MUX_2_1 . Output of 128x1 U17_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_18_output_real ;	/* Input to 2x1 U18_REAL_MUX_2_1 . Output of 128x1 U18_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_19_output_real ;	/* Input to 2x1 U19_REAL_MUX_2_1 . Output of 128x1 U19_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_20_output_real ;	/* Input to 2x1 U20_REAL_MUX_2_1 . Output of 128x1 U20_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_21_output_real ;	/* Input to 2x1 U21_REAL_MUX_2_1 . Output of 128x1 U21_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_22_output_real ;	/* Input to 2x1 U22_REAL_MUX_2_1 . Output of 128x1 U22_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_23_output_real ;	/* Input to 2x1 U23_REAL_MUX_2_1 . Output of 128x1 U23_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_24_output_real ;	/* Input to 2x1 U24_REAL_MUX_2_1 . Output of 128x1 U24_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_25_output_real ;	/* Input to 2x1 U25_REAL_MUX_2_1 . Output of 128x1 U25_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_26_output_real ;	/* Input to 2x1 U26_REAL_MUX_2_1 . Output of 128x1 U26_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_27_output_real ;	/* Input to 2x1 U27_REAL_MUX_2_1 . Output of 128x1 U27_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_28_output_real ;	/* Input to 2x1 U28_REAL_MUX_2_1 . Output of 128x1 U28_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_29_output_real ;	/* Input to 2x1 U29_REAL_MUX_2_1 . Output of 128x1 U29_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_30_output_real ;	/* Input to 2x1 U30_REAL_MUX_2_1 . Output of 128x1 U30_MUX_REAL_MEMORY */
wire [BITS-1:0] mux_31_output_real ;	/* Input to 2x1 U31_REAL_MUX_2_1 . Output of 128x1 U31_MUX_REAL_MEMORY */
wire sel_mux_2_1 ;						/* Input Selection to all insatnces of MUX_2_1 . Output of Controller  */

/*IMAG MEMORY */
/* Inputs */
wire [BITS-1:0] mux_2_1_0_output_imag ;    /* Input to Memory . Output of 2x1 U0_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_1_output_imag ;    /* Input to Memory . Output of 2x1 U1_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_2_output_imag ;    /* Input to Memory . Output of 2x1 U2_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_3_output_imag ;    /* Input to Memory . Output of 2x1 U3_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_4_output_imag ;    /* Input to Memory . Output of 2x1 U4_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_5_output_imag ;    /* Input to Memory . Output of 2x1 U5_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_6_output_imag ;    /* Input to Memory . Output of 2x1 U6_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_7_output_imag ;    /* Input to Memory . Output of 2x1 U7_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_8_output_imag ;    /* Input to Memory . Output of 2x1 U8_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_9_output_imag ;    /* Input to Memory . Output of 2x1 U9_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_10_output_imag ;    /* Input to Memory . Output of 2x1 U10_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_11_output_imag ;    /* Input to Memory . Output of 2x1 U11_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_12_output_imag ;    /* Input to Memory . Output of 2x1 U12_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_13_output_imag ;    /* Input to Memory . Output of 2x1 U13_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_14_output_imag ;    /* Input to Memory . Output of 2x1 U14_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_15_output_imag ;    /* Input to Memory . Output of 2x1 U15_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_16_output_imag ;    /* Input to Memory . Output of 2x1 U16_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_17_output_imag ;    /* Input to Memory . Output of 2x1 U17_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_18_output_imag ;    /* Input to Memory . Output of 2x1 U18_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_19_output_imag ;    /* Input to Memory . Output of 2x1 U19_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_20_output_imag ;    /* Input to Memory . Output of 2x1 U20_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_21_output_imag ;    /* Input to Memory . Output of 2x1 U21_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_22_output_imag ;    /* Input to Memory . Output of 2x1 U22_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_23_output_imag ;    /* Input to Memory . Output of 2x1 U23_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_24_output_imag ;    /* Input to Memory . Output of 2x1 U24_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_25_output_imag ;    /* Input to Memory . Output of 2x1 U25_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_26_output_imag ;    /* Input to Memory . Output of 2x1 U26_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_27_output_imag ;    /* Input to Memory . Output of 2x1 U27_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_28_output_imag ;    /* Input to Memory . Output of 2x1 U28_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_29_output_imag ;    /* Input to Memory . Output of 2x1 U29_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_30_output_imag ;    /* Input to Memory . Output of 2x1 U30_IMAG_MUX_2_1 */
wire [BITS-1:0] mux_2_1_31_output_imag ;    /* Input to Memory . Output of 2x1 U31_IMAG_MUX_2_1 */


/*Outputs*/
wire [BITS-1:0] memory_imag_output_0 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_1 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_2 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_3 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_4 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_5 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_6 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_7 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_8 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_9 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_10 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_11 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_12 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_13 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_14 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_15 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_16 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_17 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_18 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_19 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_20 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_21 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_22 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_23 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_24 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_25 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_26 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_27 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_28 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_29 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_30 ;  /* Output of Memory . Input to Registers */
wire [BITS-1:0] memory_imag_output_31 ;  /* Output of Memory . Input to Registers */


wire [BITS-1:0] mux_0_output_imag ;		/* Input to 2x1 U0_IMAG_MUX_2_1 . Output of 128x1 U0_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_1_output_imag ;		/* Input to 2x1 U1_IMAG_MUX_2_1 . Output of 128x1 U1_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_2_output_imag ;		/* Input to 2x1 U2_IMAG_MUX_2_1 . Output of 128x1 U2_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_3_output_imag ;		/* Input to 2x1 U3_IMAG_MUX_2_1 . Output of 128x1 U3_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_4_output_imag ;		/* Input to 2x1 U4_IMAG_MUX_2_1 . Output of 128x1 U4_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_5_output_imag ;		/* Input to 2x1 U5_IMAG_MUX_2_1 . Output of 128x1 U5_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_6_output_imag ;		/* Input to 2x1 U6_IMAG_MUX_2_1 . Output of 128x1 U6_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_7_output_imag ;		/* Input to 2x1 U7_IMAG_MUX_2_1 . Output of 128x1 U7_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_8_output_imag ;		/* Input to 2x1 U8_IMAG_MUX_2_1 . Output of 128x1 U8_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_9_output_imag ;		/* Input to 2x1 U9_IMAG_MUX_2_1 . Output of 128x1 U9_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_10_output_imag ;	/* Input to 2x1 U10_IMAG_MUX_2_1 . Output of 128x1 U10_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_11_output_imag ;	/* Input to 2x1 U11_IMAG_MUX_2_1 . Output of 128x1 U11_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_12_output_imag ;	/* Input to 2x1 U12_IMAG_MUX_2_1 . Output of 128x1 U12_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_13_output_imag ;	/* Input to 2x1 U13_IMAG_MUX_2_1 . Output of 128x1 U13_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_14_output_imag ;	/* Input to 2x1 U14_IMAG_MUX_2_1 . Output of 128x1 U14_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_15_output_imag ;	/* Input to 2x1 U15_IMAG_MUX_2_1 . Output of 128x1 U15_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_16_output_imag ;	/* Input to 2x1 U16_IMAG_MUX_2_1 . Output of 128x1 U16_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_17_output_imag ;	/* Input to 2x1 U17_IMAG_MUX_2_1 . Output of 128x1 U17_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_18_output_imag ;	/* Input to 2x1 U18_IMAG_MUX_2_1 . Output of 128x1 U18_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_19_output_imag ;	/* Input to 2x1 U19_IMAG_MUX_2_1 . Output of 128x1 U19_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_20_output_imag ;	/* Input to 2x1 U20_IMAG_MUX_2_1 . Output of 128x1 U20_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_21_output_imag ;	/* Input to 2x1 U21_IMAG_MUX_2_1 . Output of 128x1 U21_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_22_output_imag ;	/* Input to 2x1 U22_IMAG_MUX_2_1 . Output of 128x1 U22_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_23_output_imag ;	/* Input to 2x1 U23_IMAG_MUX_2_1 . Output of 128x1 U23_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_24_output_imag ;	/* Input to 2x1 U24_IMAG_MUX_2_1 . Output of 128x1 U24_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_25_output_imag ;	/* Input to 2x1 U25_IMAG_MUX_2_1 . Output of 128x1 U25_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_26_output_imag ;	/* Input to 2x1 U26_IMAG_MUX_2_1 . Output of 128x1 U26_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_27_output_imag ;	/* Input to 2x1 U27_IMAG_MUX_2_1 . Output of 128x1 U27_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_28_output_imag ;	/* Input to 2x1 U28_IMAG_MUX_2_1 . Output of 128x1 U28_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_29_output_imag ;	/* Input to 2x1 U29_IMAG_MUX_2_1 . Output of 128x1 U29_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_30_output_imag ;	/* Input to 2x1 U30_IMAG_MUX_2_1 . Output of 128x1 U30_MUX_IMAG_MEMORY */ 
wire [BITS-1:0] mux_31_output_imag ;	/* Input to 2x1 U31_IMAG_MUX_2_1 . Output of 128x1 U31_MUX_IMAG_MEMORY */ 



///////// output of register file . input of butterfly column//////////////
wire [BITS - 1 : 0] out_reg_r_0;
wire [BITS - 1 : 0] out_reg_r_1;
wire [BITS - 1 : 0] out_reg_r_2;
wire [BITS - 1 : 0] out_reg_r_3;
wire [BITS - 1 : 0] out_reg_r_4;
wire [BITS - 1 : 0] out_reg_r_5;
wire [BITS - 1 : 0] out_reg_r_6;
wire [BITS - 1 : 0] out_reg_r_7;
wire [BITS - 1 : 0] out_reg_r_8;
wire [BITS - 1 : 0] out_reg_r_9;
wire [BITS - 1 : 0] out_reg_r_10;
wire [BITS - 1 : 0] out_reg_r_11;
wire [BITS - 1 : 0] out_reg_r_12;
wire [BITS - 1 : 0] out_reg_r_13;
wire [BITS - 1 : 0] out_reg_r_14;
wire [BITS - 1 : 0] out_reg_r_15;
wire [BITS - 1 : 0] out_reg_r_16;
wire [BITS - 1 : 0] out_reg_r_17;
wire [BITS - 1 : 0] out_reg_r_18;
wire [BITS - 1 : 0] out_reg_r_19;
wire [BITS - 1 : 0] out_reg_r_20;
wire [BITS - 1 : 0] out_reg_r_21;
wire [BITS - 1 : 0] out_reg_r_22;
wire [BITS - 1 : 0] out_reg_r_23;
wire [BITS - 1 : 0] out_reg_r_24;
wire [BITS - 1 : 0] out_reg_r_25;
wire [BITS - 1 : 0] out_reg_r_26;
wire [BITS - 1 : 0] out_reg_r_27;
wire [BITS - 1 : 0] out_reg_r_28;
wire [BITS - 1 : 0] out_reg_r_29;
wire [BITS - 1 : 0] out_reg_r_30;
wire [BITS - 1 : 0] out_reg_r_31;
wire [BITS - 1 : 0] out_reg_r_32;
wire [BITS - 1 : 0] out_reg_r_33;
wire [BITS - 1 : 0] out_reg_r_34;
wire [BITS - 1 : 0] out_reg_r_35;
wire [BITS - 1 : 0] out_reg_r_36;
wire [BITS - 1 : 0] out_reg_r_37;
wire [BITS - 1 : 0] out_reg_r_38;
wire [BITS - 1 : 0] out_reg_r_39;
wire [BITS - 1 : 0] out_reg_r_40;
wire [BITS - 1 : 0] out_reg_r_41;
wire [BITS - 1 : 0] out_reg_r_42;
wire [BITS - 1 : 0] out_reg_r_43;
wire [BITS - 1 : 0] out_reg_r_44;
wire [BITS - 1 : 0] out_reg_r_45;
wire [BITS - 1 : 0] out_reg_r_46;
wire [BITS - 1 : 0] out_reg_r_47;
wire [BITS - 1 : 0] out_reg_r_48;
wire [BITS - 1 : 0] out_reg_r_49;
wire [BITS - 1 : 0] out_reg_r_50;
wire [BITS - 1 : 0] out_reg_r_51;
wire [BITS - 1 : 0] out_reg_r_52;
wire [BITS - 1 : 0] out_reg_r_53;
wire [BITS - 1 : 0] out_reg_r_54;
wire [BITS - 1 : 0] out_reg_r_55;
wire [BITS - 1 : 0] out_reg_r_56;
wire [BITS - 1 : 0] out_reg_r_57;
wire [BITS - 1 : 0] out_reg_r_58;
wire [BITS - 1 : 0] out_reg_r_59;
wire [BITS - 1 : 0] out_reg_r_60;
wire [BITS - 1 : 0] out_reg_r_61;
wire [BITS - 1 : 0] out_reg_r_62;
wire [BITS - 1 : 0] out_reg_r_63;
wire [BITS - 1 : 0] out_reg_r_64;
wire [BITS - 1 : 0] out_reg_r_65;
wire [BITS - 1 : 0] out_reg_r_66;
wire [BITS - 1 : 0] out_reg_r_67;
wire [BITS - 1 : 0] out_reg_r_68;
wire [BITS - 1 : 0] out_reg_r_69;
wire [BITS - 1 : 0] out_reg_r_70;
wire [BITS - 1 : 0] out_reg_r_71;
wire [BITS - 1 : 0] out_reg_r_72;
wire [BITS - 1 : 0] out_reg_r_73;
wire [BITS - 1 : 0] out_reg_r_74;
wire [BITS - 1 : 0] out_reg_r_75;
wire [BITS - 1 : 0] out_reg_r_76;
wire [BITS - 1 : 0] out_reg_r_77;
wire [BITS - 1 : 0] out_reg_r_78;
wire [BITS - 1 : 0] out_reg_r_79;
wire [BITS - 1 : 0] out_reg_r_80;
wire [BITS - 1 : 0] out_reg_r_81;
wire [BITS - 1 : 0] out_reg_r_82;
wire [BITS - 1 : 0] out_reg_r_83;
wire [BITS - 1 : 0] out_reg_r_84;
wire [BITS - 1 : 0] out_reg_r_85;
wire [BITS - 1 : 0] out_reg_r_86;
wire [BITS - 1 : 0] out_reg_r_87;
wire [BITS - 1 : 0] out_reg_r_88;
wire [BITS - 1 : 0] out_reg_r_89;
wire [BITS - 1 : 0] out_reg_r_90;
wire [BITS - 1 : 0] out_reg_r_91;
wire [BITS - 1 : 0] out_reg_r_92;
wire [BITS - 1 : 0] out_reg_r_93;
wire [BITS - 1 : 0] out_reg_r_94;
wire [BITS - 1 : 0] out_reg_r_95;
wire [BITS - 1 : 0] out_reg_r_96;
wire [BITS - 1 : 0] out_reg_r_97;
wire [BITS - 1 : 0] out_reg_r_98;
wire [BITS - 1 : 0] out_reg_r_99;
wire [BITS - 1 : 0] out_reg_r_100;
wire [BITS - 1 : 0] out_reg_r_101;
wire [BITS - 1 : 0] out_reg_r_102;
wire [BITS - 1 : 0] out_reg_r_103;
wire [BITS - 1 : 0] out_reg_r_104;
wire [BITS - 1 : 0] out_reg_r_105;
wire [BITS - 1 : 0] out_reg_r_106;
wire [BITS - 1 : 0] out_reg_r_107;
wire [BITS - 1 : 0] out_reg_r_108;
wire [BITS - 1 : 0] out_reg_r_109;
wire [BITS - 1 : 0] out_reg_r_110;
wire [BITS - 1 : 0] out_reg_r_111;
wire [BITS - 1 : 0] out_reg_r_112;
wire [BITS - 1 : 0] out_reg_r_113;
wire [BITS - 1 : 0] out_reg_r_114;
wire [BITS - 1 : 0] out_reg_r_115;
wire [BITS - 1 : 0] out_reg_r_116;
wire [BITS - 1 : 0] out_reg_r_117;
wire [BITS - 1 : 0] out_reg_r_118;
wire [BITS - 1 : 0] out_reg_r_119;
wire [BITS - 1 : 0] out_reg_r_120;
wire [BITS - 1 : 0] out_reg_r_121;
wire [BITS - 1 : 0] out_reg_r_122;
wire [BITS - 1 : 0] out_reg_r_123;
wire [BITS - 1 : 0] out_reg_r_124;
wire [BITS - 1 : 0] out_reg_r_125;
wire [BITS - 1 : 0] out_reg_r_126;
wire [BITS - 1 : 0] out_reg_r_127;


wire [BITS - 1 : 0] out_reg_i_0;		/*Output of Register File and Input to Butterfly Column Top */
wire [BITS - 1 : 0] out_reg_i_1;
wire [BITS - 1 : 0] out_reg_i_2;
wire [BITS - 1 : 0] out_reg_i_3;
wire [BITS - 1 : 0] out_reg_i_4;
wire [BITS - 1 : 0] out_reg_i_5;
wire [BITS - 1 : 0] out_reg_i_6;
wire [BITS - 1 : 0] out_reg_i_7;
wire [BITS - 1 : 0] out_reg_i_8;
wire [BITS - 1 : 0] out_reg_i_9;
wire [BITS - 1 : 0] out_reg_i_10;
wire [BITS - 1 : 0] out_reg_i_11;
wire [BITS - 1 : 0] out_reg_i_12;
wire [BITS - 1 : 0] out_reg_i_13;
wire [BITS - 1 : 0] out_reg_i_14;
wire [BITS - 1 : 0] out_reg_i_15;
wire [BITS - 1 : 0] out_reg_i_16;
wire [BITS - 1 : 0] out_reg_i_17;
wire [BITS - 1 : 0] out_reg_i_18;
wire [BITS - 1 : 0] out_reg_i_19;
wire [BITS - 1 : 0] out_reg_i_20;
wire [BITS - 1 : 0] out_reg_i_21;
wire [BITS - 1 : 0] out_reg_i_22;
wire [BITS - 1 : 0] out_reg_i_23;
wire [BITS - 1 : 0] out_reg_i_24;
wire [BITS - 1 : 0] out_reg_i_25;
wire [BITS - 1 : 0] out_reg_i_26;
wire [BITS - 1 : 0] out_reg_i_27;
wire [BITS - 1 : 0] out_reg_i_28;
wire [BITS - 1 : 0] out_reg_i_29;
wire [BITS - 1 : 0] out_reg_i_30;
wire [BITS - 1 : 0] out_reg_i_31;
wire [BITS - 1 : 0] out_reg_i_32;
wire [BITS - 1 : 0] out_reg_i_33;
wire [BITS - 1 : 0] out_reg_i_34;
wire [BITS - 1 : 0] out_reg_i_35;
wire [BITS - 1 : 0] out_reg_i_36;
wire [BITS - 1 : 0] out_reg_i_37;
wire [BITS - 1 : 0] out_reg_i_38;
wire [BITS - 1 : 0] out_reg_i_39;
wire [BITS - 1 : 0] out_reg_i_40;
wire [BITS - 1 : 0] out_reg_i_41;
wire [BITS - 1 : 0] out_reg_i_42;
wire [BITS - 1 : 0] out_reg_i_43;
wire [BITS - 1 : 0] out_reg_i_44;
wire [BITS - 1 : 0] out_reg_i_45;
wire [BITS - 1 : 0] out_reg_i_46;
wire [BITS - 1 : 0] out_reg_i_47;
wire [BITS - 1 : 0] out_reg_i_48;
wire [BITS - 1 : 0] out_reg_i_49;
wire [BITS - 1 : 0] out_reg_i_50;
wire [BITS - 1 : 0] out_reg_i_51;
wire [BITS - 1 : 0] out_reg_i_52;
wire [BITS - 1 : 0] out_reg_i_53;
wire [BITS - 1 : 0] out_reg_i_54;
wire [BITS - 1 : 0] out_reg_i_55;
wire [BITS - 1 : 0] out_reg_i_56;
wire [BITS - 1 : 0] out_reg_i_57;
wire [BITS - 1 : 0] out_reg_i_58;
wire [BITS - 1 : 0] out_reg_i_59;
wire [BITS - 1 : 0] out_reg_i_60;
wire [BITS - 1 : 0] out_reg_i_61;
wire [BITS - 1 : 0] out_reg_i_62;
wire [BITS - 1 : 0] out_reg_i_63;
wire [BITS - 1 : 0] out_reg_i_64;
wire [BITS - 1 : 0] out_reg_i_65;
wire [BITS - 1 : 0] out_reg_i_66;
wire [BITS - 1 : 0] out_reg_i_67;
wire [BITS - 1 : 0] out_reg_i_68;
wire [BITS - 1 : 0] out_reg_i_69;
wire [BITS - 1 : 0] out_reg_i_70;
wire [BITS - 1 : 0] out_reg_i_71;
wire [BITS - 1 : 0] out_reg_i_72;
wire [BITS - 1 : 0] out_reg_i_73;
wire [BITS - 1 : 0] out_reg_i_74;
wire [BITS - 1 : 0] out_reg_i_75;
wire [BITS - 1 : 0] out_reg_i_76;
wire [BITS - 1 : 0] out_reg_i_77;
wire [BITS - 1 : 0] out_reg_i_78;
wire [BITS - 1 : 0] out_reg_i_79;
wire [BITS - 1 : 0] out_reg_i_80;
wire [BITS - 1 : 0] out_reg_i_81;
wire [BITS - 1 : 0] out_reg_i_82;
wire [BITS - 1 : 0] out_reg_i_83;
wire [BITS - 1 : 0] out_reg_i_84;
wire [BITS - 1 : 0] out_reg_i_85;
wire [BITS - 1 : 0] out_reg_i_86;
wire [BITS - 1 : 0] out_reg_i_87;
wire [BITS - 1 : 0] out_reg_i_88;
wire [BITS - 1 : 0] out_reg_i_89;
wire [BITS - 1 : 0] out_reg_i_90;
wire [BITS - 1 : 0] out_reg_i_91;
wire [BITS - 1 : 0] out_reg_i_92;
wire [BITS - 1 : 0] out_reg_i_93;
wire [BITS - 1 : 0] out_reg_i_94;
wire [BITS - 1 : 0] out_reg_i_95;
wire [BITS - 1 : 0] out_reg_i_96;
wire [BITS - 1 : 0] out_reg_i_97;
wire [BITS - 1 : 0] out_reg_i_98;
wire [BITS - 1 : 0] out_reg_i_99;
wire [BITS - 1 : 0] out_reg_i_100;
wire [BITS - 1 : 0] out_reg_i_101;
wire [BITS - 1 : 0] out_reg_i_102;
wire [BITS - 1 : 0] out_reg_i_103;
wire [BITS - 1 : 0] out_reg_i_104;
wire [BITS - 1 : 0] out_reg_i_105;
wire [BITS - 1 : 0] out_reg_i_106;
wire [BITS - 1 : 0] out_reg_i_107;
wire [BITS - 1 : 0] out_reg_i_108;
wire [BITS - 1 : 0] out_reg_i_109;
wire [BITS - 1 : 0] out_reg_i_110;
wire [BITS - 1 : 0] out_reg_i_111;
wire [BITS - 1 : 0] out_reg_i_112;
wire [BITS - 1 : 0] out_reg_i_113;
wire [BITS - 1 : 0] out_reg_i_114;
wire [BITS - 1 : 0] out_reg_i_115;
wire [BITS - 1 : 0] out_reg_i_116;
wire [BITS - 1 : 0] out_reg_i_117;
wire [BITS - 1 : 0] out_reg_i_118;
wire [BITS - 1 : 0] out_reg_i_119;
wire [BITS - 1 : 0] out_reg_i_120;
wire [BITS - 1 : 0] out_reg_i_121;
wire [BITS - 1 : 0] out_reg_i_122;
wire [BITS - 1 : 0] out_reg_i_123;
wire [BITS - 1 : 0] out_reg_i_124;
wire [BITS - 1 : 0] out_reg_i_125;
wire [BITS - 1 : 0] out_reg_i_126;
wire [BITS - 1 : 0] out_reg_i_127;



////output of twiddle register . input of butterfly column
wire [BITS - 1 : 0] out_reg_twiddle_r_0;
wire [BITS - 1 : 0] out_reg_twiddle_i_0;
wire [BITS - 1 : 0] out_reg_twiddle_r_1;
wire [BITS - 1 : 0] out_reg_twiddle_i_1;
wire [BITS - 1 : 0] out_reg_twiddle_r_2;
wire [BITS - 1 : 0] out_reg_twiddle_i_2;
wire [BITS - 1 : 0] out_reg_twiddle_r_3;
wire [BITS - 1 : 0] out_reg_twiddle_i_3;
wire [BITS - 1 : 0] out_reg_twiddle_r_4;
wire [BITS - 1 : 0] out_reg_twiddle_i_4;
wire [BITS - 1 : 0] out_reg_twiddle_r_5;
wire [BITS - 1 : 0] out_reg_twiddle_i_5;
wire [BITS - 1 : 0] out_reg_twiddle_r_6;
wire [BITS - 1 : 0] out_reg_twiddle_i_6;
wire [BITS - 1 : 0] out_reg_twiddle_r_7;
wire [BITS - 1 : 0] out_reg_twiddle_i_7;
wire [BITS - 1 : 0] out_reg_twiddle_r_8;
wire [BITS - 1 : 0] out_reg_twiddle_i_8;
wire [BITS - 1 : 0] out_reg_twiddle_r_9;
wire [BITS - 1 : 0] out_reg_twiddle_i_9;
wire [BITS - 1 : 0] out_reg_twiddle_r_10;
wire [BITS - 1 : 0] out_reg_twiddle_i_10;
wire [BITS - 1 : 0] out_reg_twiddle_r_11;
wire [BITS - 1 : 0] out_reg_twiddle_i_11;
wire [BITS - 1 : 0] out_reg_twiddle_r_12;
wire [BITS - 1 : 0] out_reg_twiddle_i_12;
wire [BITS - 1 : 0] out_reg_twiddle_r_13;
wire [BITS - 1 : 0] out_reg_twiddle_i_13;
wire [BITS - 1 : 0] out_reg_twiddle_r_14;
wire [BITS - 1 : 0] out_reg_twiddle_i_14;
wire [BITS - 1 : 0] out_reg_twiddle_r_15;
wire [BITS - 1 : 0] out_reg_twiddle_i_15;
wire [BITS - 1 : 0] out_reg_twiddle_r_16;
wire [BITS - 1 : 0] out_reg_twiddle_i_16;
wire [BITS - 1 : 0] out_reg_twiddle_r_17;
wire [BITS - 1 : 0] out_reg_twiddle_i_17;
wire [BITS - 1 : 0] out_reg_twiddle_r_18;
wire [BITS - 1 : 0] out_reg_twiddle_i_18;
wire [BITS - 1 : 0] out_reg_twiddle_r_19;
wire [BITS - 1 : 0] out_reg_twiddle_i_19;
wire [BITS - 1 : 0] out_reg_twiddle_r_20;
wire [BITS - 1 : 0] out_reg_twiddle_i_20;
wire [BITS - 1 : 0] out_reg_twiddle_r_21;
wire [BITS - 1 : 0] out_reg_twiddle_i_21;
wire [BITS - 1 : 0] out_reg_twiddle_r_22;
wire [BITS - 1 : 0] out_reg_twiddle_i_22;
wire [BITS - 1 : 0] out_reg_twiddle_r_23;
wire [BITS - 1 : 0] out_reg_twiddle_i_23;
wire [BITS - 1 : 0] out_reg_twiddle_r_24;
wire [BITS - 1 : 0] out_reg_twiddle_i_24;
wire [BITS - 1 : 0] out_reg_twiddle_r_25;
wire [BITS - 1 : 0] out_reg_twiddle_i_25;
wire [BITS - 1 : 0] out_reg_twiddle_r_26;
wire [BITS - 1 : 0] out_reg_twiddle_i_26;
wire [BITS - 1 : 0] out_reg_twiddle_r_27;
wire [BITS - 1 : 0] out_reg_twiddle_i_27;
wire [BITS - 1 : 0] out_reg_twiddle_r_28;
wire [BITS - 1 : 0] out_reg_twiddle_i_28;
wire [BITS - 1 : 0] out_reg_twiddle_r_29;
wire [BITS - 1 : 0] out_reg_twiddle_i_29;
wire [BITS - 1 : 0] out_reg_twiddle_r_30;
wire [BITS - 1 : 0] out_reg_twiddle_i_30;
wire [BITS - 1 : 0] out_reg_twiddle_r_31;
wire [BITS - 1 : 0] out_reg_twiddle_i_31;
wire [BITS - 1 : 0] out_reg_twiddle_r_32;
wire [BITS - 1 : 0] out_reg_twiddle_i_32;
wire [BITS - 1 : 0] out_reg_twiddle_r_33;
wire [BITS - 1 : 0] out_reg_twiddle_i_33;
wire [BITS - 1 : 0] out_reg_twiddle_r_34;
wire [BITS - 1 : 0] out_reg_twiddle_i_34;
wire [BITS - 1 : 0] out_reg_twiddle_r_35;
wire [BITS - 1 : 0] out_reg_twiddle_i_35;
wire [BITS - 1 : 0] out_reg_twiddle_r_36;
wire [BITS - 1 : 0] out_reg_twiddle_i_36;
wire [BITS - 1 : 0] out_reg_twiddle_r_37;
wire [BITS - 1 : 0] out_reg_twiddle_i_37;
wire [BITS - 1 : 0] out_reg_twiddle_r_38;
wire [BITS - 1 : 0] out_reg_twiddle_i_38;
wire [BITS - 1 : 0] out_reg_twiddle_r_39;
wire [BITS - 1 : 0] out_reg_twiddle_i_39;
wire [BITS - 1 : 0] out_reg_twiddle_r_40;
wire [BITS - 1 : 0] out_reg_twiddle_i_40;
wire [BITS - 1 : 0] out_reg_twiddle_r_41;
wire [BITS - 1 : 0] out_reg_twiddle_i_41;
wire [BITS - 1 : 0] out_reg_twiddle_r_42;
wire [BITS - 1 : 0] out_reg_twiddle_i_42;
wire [BITS - 1 : 0] out_reg_twiddle_r_43;
wire [BITS - 1 : 0] out_reg_twiddle_i_43;
wire [BITS - 1 : 0] out_reg_twiddle_r_44;
wire [BITS - 1 : 0] out_reg_twiddle_i_44;
wire [BITS - 1 : 0] out_reg_twiddle_r_45;
wire [BITS - 1 : 0] out_reg_twiddle_i_45;
wire [BITS - 1 : 0] out_reg_twiddle_r_46;
wire [BITS - 1 : 0] out_reg_twiddle_i_46;
wire [BITS - 1 : 0] out_reg_twiddle_r_47;
wire [BITS - 1 : 0] out_reg_twiddle_i_47;
wire [BITS - 1 : 0] out_reg_twiddle_r_48;
wire [BITS - 1 : 0] out_reg_twiddle_i_48;
wire [BITS - 1 : 0] out_reg_twiddle_r_49;
wire [BITS - 1 : 0] out_reg_twiddle_i_49;
wire [BITS - 1 : 0] out_reg_twiddle_r_50;
wire [BITS - 1 : 0] out_reg_twiddle_i_50;
wire [BITS - 1 : 0] out_reg_twiddle_r_51;
wire [BITS - 1 : 0] out_reg_twiddle_i_51;
wire [BITS - 1 : 0] out_reg_twiddle_r_52;
wire [BITS - 1 : 0] out_reg_twiddle_i_52;
wire [BITS - 1 : 0] out_reg_twiddle_r_53;
wire [BITS - 1 : 0] out_reg_twiddle_i_53;
wire [BITS - 1 : 0] out_reg_twiddle_r_54;
wire [BITS - 1 : 0] out_reg_twiddle_i_54;
wire [BITS - 1 : 0] out_reg_twiddle_r_55;
wire [BITS - 1 : 0] out_reg_twiddle_i_55;
wire [BITS - 1 : 0] out_reg_twiddle_r_56;
wire [BITS - 1 : 0] out_reg_twiddle_i_56;
wire [BITS - 1 : 0] out_reg_twiddle_r_57;
wire [BITS - 1 : 0] out_reg_twiddle_i_57;
wire [BITS - 1 : 0] out_reg_twiddle_r_58;
wire [BITS - 1 : 0] out_reg_twiddle_i_58;
wire [BITS - 1 : 0] out_reg_twiddle_r_59;
wire [BITS - 1 : 0] out_reg_twiddle_i_59;
wire [BITS - 1 : 0] out_reg_twiddle_r_60;
wire [BITS - 1 : 0] out_reg_twiddle_i_60;
wire [BITS - 1 : 0] out_reg_twiddle_r_61;
wire [BITS - 1 : 0] out_reg_twiddle_i_61;
wire [BITS - 1 : 0] out_reg_twiddle_r_62;
wire [BITS - 1 : 0] out_reg_twiddle_i_62;
wire [BITS - 1 : 0] out_reg_twiddle_r_63;
wire [BITS - 1 : 0] out_reg_twiddle_i_63;


////output of twiddle ROM . input of twiddle register

wire [BITS - 1 : 0] ROM_out_twiddle_r_0;
wire [BITS - 1 : 0] ROM_out_twiddle_i_0;
wire [BITS - 1 : 0] ROM_out_twiddle_r_1;
wire [BITS - 1 : 0] ROM_out_twiddle_i_1;
wire [BITS - 1 : 0] ROM_out_twiddle_r_2;
wire [BITS - 1 : 0] ROM_out_twiddle_i_2;
wire [BITS - 1 : 0] ROM_out_twiddle_r_3;
wire [BITS - 1 : 0] ROM_out_twiddle_i_3;
wire [BITS - 1 : 0] ROM_out_twiddle_r_4;
wire [BITS - 1 : 0] ROM_out_twiddle_i_4;
wire [BITS - 1 : 0] ROM_out_twiddle_r_5;
wire [BITS - 1 : 0] ROM_out_twiddle_i_5;
wire [BITS - 1 : 0] ROM_out_twiddle_r_6;
wire [BITS - 1 : 0] ROM_out_twiddle_i_6;
wire [BITS - 1 : 0] ROM_out_twiddle_r_7;
wire [BITS - 1 : 0] ROM_out_twiddle_i_7;
wire [BITS - 1 : 0] ROM_out_twiddle_r_8;
wire [BITS - 1 : 0] ROM_out_twiddle_i_8;
wire [BITS - 1 : 0] ROM_out_twiddle_r_9;
wire [BITS - 1 : 0] ROM_out_twiddle_i_9;
wire [BITS - 1 : 0] ROM_out_twiddle_r_10;
wire [BITS - 1 : 0] ROM_out_twiddle_i_10;
wire [BITS - 1 : 0] ROM_out_twiddle_r_11;
wire [BITS - 1 : 0] ROM_out_twiddle_i_11;
wire [BITS - 1 : 0] ROM_out_twiddle_r_12;
wire [BITS - 1 : 0] ROM_out_twiddle_i_12;
wire [BITS - 1 : 0] ROM_out_twiddle_r_13;
wire [BITS - 1 : 0] ROM_out_twiddle_i_13;
wire [BITS - 1 : 0] ROM_out_twiddle_r_14;
wire [BITS - 1 : 0] ROM_out_twiddle_i_14;
wire [BITS - 1 : 0] ROM_out_twiddle_r_15;
wire [BITS - 1 : 0] ROM_out_twiddle_i_15;


//MUX_4_1 output . MUX_2_1 input

wire [BITS - 1 : 0] mux4_mux2_0_r;		/* Inputs to 2x1 MUX. Outputs of 4x1 MUX */
wire [BITS - 1 : 0] mux4_mux2_0_i;
wire [BITS - 1 : 0] mux4_mux2_1_r;
wire [BITS - 1 : 0] mux4_mux2_1_i;
wire [BITS - 1 : 0] mux4_mux2_2_r;
wire [BITS - 1 : 0] mux4_mux2_2_i;
wire [BITS - 1 : 0] mux4_mux2_3_r;
wire [BITS - 1 : 0] mux4_mux2_3_i;
wire [BITS - 1 : 0] mux4_mux2_4_r;
wire [BITS - 1 : 0] mux4_mux2_4_i;
wire [BITS - 1 : 0] mux4_mux2_5_r;
wire [BITS - 1 : 0] mux4_mux2_5_i;
wire [BITS - 1 : 0] mux4_mux2_6_r;
wire [BITS - 1 : 0] mux4_mux2_6_i;
wire [BITS - 1 : 0] mux4_mux2_7_r;
wire [BITS - 1 : 0] mux4_mux2_7_i;
wire [BITS - 1 : 0] mux4_mux2_8_r;
wire [BITS - 1 : 0] mux4_mux2_8_i;
wire [BITS - 1 : 0] mux4_mux2_9_r;
wire [BITS - 1 : 0] mux4_mux2_9_i;
wire [BITS - 1 : 0] mux4_mux2_10_r;
wire [BITS - 1 : 0] mux4_mux2_10_i;
wire [BITS - 1 : 0] mux4_mux2_11_r;
wire [BITS - 1 : 0] mux4_mux2_11_i;
wire [BITS - 1 : 0] mux4_mux2_12_r;
wire [BITS - 1 : 0] mux4_mux2_12_i;
wire [BITS - 1 : 0] mux4_mux2_13_r;
wire [BITS - 1 : 0] mux4_mux2_13_i;
wire [BITS - 1 : 0] mux4_mux2_14_r;
wire [BITS - 1 : 0] mux4_mux2_14_i;
wire [BITS - 1 : 0] mux4_mux2_15_r;
wire [BITS - 1 : 0] mux4_mux2_15_i;
wire [BITS - 1 : 0] mux4_mux2_16_r;
wire [BITS - 1 : 0] mux4_mux2_16_i;
wire [BITS - 1 : 0] mux4_mux2_17_r;
wire [BITS - 1 : 0] mux4_mux2_17_i;
wire [BITS - 1 : 0] mux4_mux2_18_r;
wire [BITS - 1 : 0] mux4_mux2_18_i;
wire [BITS - 1 : 0] mux4_mux2_19_r;
wire [BITS - 1 : 0] mux4_mux2_19_i;
wire [BITS - 1 : 0] mux4_mux2_20_r;
wire [BITS - 1 : 0] mux4_mux2_20_i;
wire [BITS - 1 : 0] mux4_mux2_21_r;
wire [BITS - 1 : 0] mux4_mux2_21_i;
wire [BITS - 1 : 0] mux4_mux2_22_r;
wire [BITS - 1 : 0] mux4_mux2_22_i;
wire [BITS - 1 : 0] mux4_mux2_23_r;
wire [BITS - 1 : 0] mux4_mux2_23_i;
wire [BITS - 1 : 0] mux4_mux2_24_r;
wire [BITS - 1 : 0] mux4_mux2_24_i;
wire [BITS - 1 : 0] mux4_mux2_25_r;
wire [BITS - 1 : 0] mux4_mux2_25_i;
wire [BITS - 1 : 0] mux4_mux2_26_r;
wire [BITS - 1 : 0] mux4_mux2_26_i;
wire [BITS - 1 : 0] mux4_mux2_27_r;
wire [BITS - 1 : 0] mux4_mux2_27_i;
wire [BITS - 1 : 0] mux4_mux2_28_r;
wire [BITS - 1 : 0] mux4_mux2_28_i;
wire [BITS - 1 : 0] mux4_mux2_29_r;
wire [BITS - 1 : 0] mux4_mux2_29_i;
wire [BITS - 1 : 0] mux4_mux2_30_r;
wire [BITS - 1 : 0] mux4_mux2_30_i;
wire [BITS - 1 : 0] mux4_mux2_31_r;
wire [BITS - 1 : 0] mux4_mux2_31_i;


  




Reg_File #(.BITS(BITS),.NUMBER_OF_REGISTERS(NUMBER_OF_ENABLE_BITS)) Reg_File_REAL 
( 

.WrEn(reg_en) , 
.clk(clk) ,
.rst(rst) , 
  
.WrData_0(memory_real_output_0),
.WrData_1(memory_real_output_0),
.WrData_2(memory_real_output_0),
.WrData_3(memory_real_output_0),
.WrData_4(memory_real_output_1),
.WrData_5(memory_real_output_1),
.WrData_6(memory_real_output_1),
.WrData_7(memory_real_output_1),
.WrData_8(memory_real_output_2),
.WrData_9(memory_real_output_2),
.WrData_10(memory_real_output_2),
.WrData_11(memory_real_output_2),
.WrData_12(memory_real_output_3),
.WrData_13(memory_real_output_3),
.WrData_14(memory_real_output_3),
.WrData_15(memory_real_output_3),
.WrData_16(memory_real_output_4),
.WrData_17(memory_real_output_4),
.WrData_18(memory_real_output_4),
.WrData_19(memory_real_output_4),
.WrData_20(memory_real_output_5),
.WrData_21(memory_real_output_5),
.WrData_22(memory_real_output_5),
.WrData_23(memory_real_output_5),
.WrData_24(memory_real_output_6),
.WrData_25(memory_real_output_6),
.WrData_26(memory_real_output_6),
.WrData_27(memory_real_output_6),
.WrData_28(memory_real_output_7),
.WrData_29(memory_real_output_7),
.WrData_30(memory_real_output_7),
.WrData_31(memory_real_output_7),
.WrData_32(memory_real_output_8),
.WrData_33(memory_real_output_8),
.WrData_34(memory_real_output_8),
.WrData_35(memory_real_output_8),
.WrData_36(memory_real_output_9),
.WrData_37(memory_real_output_9),
.WrData_38(memory_real_output_9),
.WrData_39(memory_real_output_9),
.WrData_40(memory_real_output_10),
.WrData_41(memory_real_output_10),
.WrData_42(memory_real_output_10),
.WrData_43(memory_real_output_10),
.WrData_44(memory_real_output_11),
.WrData_45(memory_real_output_11),
.WrData_46(memory_real_output_11),
.WrData_47(memory_real_output_11),
.WrData_48(memory_real_output_12),
.WrData_49(memory_real_output_12),
.WrData_50(memory_real_output_12),
.WrData_51(memory_real_output_12),
.WrData_52(memory_real_output_13),
.WrData_53(memory_real_output_13),
.WrData_54(memory_real_output_13),
.WrData_55(memory_real_output_13),
.WrData_56(memory_real_output_14),
.WrData_57(memory_real_output_14),
.WrData_58(memory_real_output_14),
.WrData_59(memory_real_output_14),
.WrData_60(memory_real_output_15),
.WrData_61(memory_real_output_15),
.WrData_62(memory_real_output_15),
.WrData_63(memory_real_output_15),
.WrData_64(memory_real_output_16),
.WrData_65(memory_real_output_16),
.WrData_66(memory_real_output_16),
.WrData_67(memory_real_output_16),
.WrData_68(memory_real_output_17),
.WrData_69(memory_real_output_17),
.WrData_70(memory_real_output_17),
.WrData_71(memory_real_output_17),
.WrData_72(memory_real_output_18),
.WrData_73(memory_real_output_18),
.WrData_74(memory_real_output_18),
.WrData_75(memory_real_output_18),
.WrData_76(memory_real_output_19),
.WrData_77(memory_real_output_19),
.WrData_78(memory_real_output_19),
.WrData_79(memory_real_output_19),
.WrData_80(memory_real_output_20),
.WrData_81(memory_real_output_20),
.WrData_82(memory_real_output_20),
.WrData_83(memory_real_output_20),
.WrData_84(memory_real_output_21),
.WrData_85(memory_real_output_21),
.WrData_86(memory_real_output_21),
.WrData_87(memory_real_output_21),
.WrData_88(memory_real_output_22),
.WrData_89(memory_real_output_22),
.WrData_90(memory_real_output_22),
.WrData_91(memory_real_output_22),
.WrData_92(memory_real_output_23),
.WrData_93(memory_real_output_23),
.WrData_94(memory_real_output_23),
.WrData_95(memory_real_output_23),
.WrData_96(memory_real_output_24),
.WrData_97(memory_real_output_24),
.WrData_98(memory_real_output_24),
.WrData_99(memory_real_output_24),
.WrData_100(memory_real_output_25),
.WrData_101(memory_real_output_25),
.WrData_102(memory_real_output_25),
.WrData_103(memory_real_output_25),
.WrData_104(memory_real_output_26),
.WrData_105(memory_real_output_26),
.WrData_106(memory_real_output_26),
.WrData_107(memory_real_output_26),
.WrData_108(memory_real_output_27),
.WrData_109(memory_real_output_27),
.WrData_110(memory_real_output_27),
.WrData_111(memory_real_output_27),
.WrData_112(memory_real_output_28),
.WrData_113(memory_real_output_28),
.WrData_114(memory_real_output_28),
.WrData_115(memory_real_output_28),
.WrData_116(memory_real_output_29),
.WrData_117(memory_real_output_29),
.WrData_118(memory_real_output_29),
.WrData_119(memory_real_output_29),
.WrData_120(memory_real_output_30),
.WrData_121(memory_real_output_30),
.WrData_122(memory_real_output_30),
.WrData_123(memory_real_output_30),
.WrData_124(memory_real_output_31),
.WrData_125(memory_real_output_31),
.WrData_126(memory_real_output_31),
.WrData_127(memory_real_output_31),


.RdData_0(out_reg_r_0),
.RdData_1(out_reg_r_1),
.RdData_2(out_reg_r_2),
.RdData_3(out_reg_r_3),
.RdData_4(out_reg_r_4),
.RdData_5(out_reg_r_5),
.RdData_6(out_reg_r_6),
.RdData_7(out_reg_r_7),
.RdData_8(out_reg_r_8),
.RdData_9(out_reg_r_9),
.RdData_10(out_reg_r_10),
.RdData_11(out_reg_r_11),
.RdData_12(out_reg_r_12),
.RdData_13(out_reg_r_13),
.RdData_14(out_reg_r_14),
.RdData_15(out_reg_r_15),
.RdData_16(out_reg_r_16),
.RdData_17(out_reg_r_17),
.RdData_18(out_reg_r_18),
.RdData_19(out_reg_r_19),
.RdData_20(out_reg_r_20),
.RdData_21(out_reg_r_21),
.RdData_22(out_reg_r_22),
.RdData_23(out_reg_r_23),
.RdData_24(out_reg_r_24),
.RdData_25(out_reg_r_25),
.RdData_26(out_reg_r_26),
.RdData_27(out_reg_r_27),
.RdData_28(out_reg_r_28),
.RdData_29(out_reg_r_29),
.RdData_30(out_reg_r_30),
.RdData_31(out_reg_r_31),
.RdData_32(out_reg_r_32),
.RdData_33(out_reg_r_33),
.RdData_34(out_reg_r_34),
.RdData_35(out_reg_r_35),
.RdData_36(out_reg_r_36),
.RdData_37(out_reg_r_37),
.RdData_38(out_reg_r_38),
.RdData_39(out_reg_r_39),
.RdData_40(out_reg_r_40),
.RdData_41(out_reg_r_41),
.RdData_42(out_reg_r_42),
.RdData_43(out_reg_r_43),
.RdData_44(out_reg_r_44),
.RdData_45(out_reg_r_45),
.RdData_46(out_reg_r_46),
.RdData_47(out_reg_r_47),
.RdData_48(out_reg_r_48),
.RdData_49(out_reg_r_49),
.RdData_50(out_reg_r_50),
.RdData_51(out_reg_r_51),
.RdData_52(out_reg_r_52),
.RdData_53(out_reg_r_53),
.RdData_54(out_reg_r_54),
.RdData_55(out_reg_r_55),
.RdData_56(out_reg_r_56),
.RdData_57(out_reg_r_57),
.RdData_58(out_reg_r_58),
.RdData_59(out_reg_r_59),
.RdData_60(out_reg_r_60),
.RdData_61(out_reg_r_61),
.RdData_62(out_reg_r_62),
.RdData_63(out_reg_r_63),
.RdData_64(out_reg_r_64),
.RdData_65(out_reg_r_65),
.RdData_66(out_reg_r_66),
.RdData_67(out_reg_r_67),
.RdData_68(out_reg_r_68),
.RdData_69(out_reg_r_69),
.RdData_70(out_reg_r_70),
.RdData_71(out_reg_r_71),
.RdData_72(out_reg_r_72),
.RdData_73(out_reg_r_73),
.RdData_74(out_reg_r_74),
.RdData_75(out_reg_r_75),
.RdData_76(out_reg_r_76),
.RdData_77(out_reg_r_77),
.RdData_78(out_reg_r_78),
.RdData_79(out_reg_r_79),
.RdData_80(out_reg_r_80),
.RdData_81(out_reg_r_81),
.RdData_82(out_reg_r_82),
.RdData_83(out_reg_r_83),
.RdData_84(out_reg_r_84),
.RdData_85(out_reg_r_85),
.RdData_86(out_reg_r_86),
.RdData_87(out_reg_r_87),
.RdData_88(out_reg_r_88),
.RdData_89(out_reg_r_89),
.RdData_90(out_reg_r_90),
.RdData_91(out_reg_r_91),
.RdData_92(out_reg_r_92),
.RdData_93(out_reg_r_93),
.RdData_94(out_reg_r_94),
.RdData_95(out_reg_r_95),
.RdData_96(out_reg_r_96),
.RdData_97(out_reg_r_97),
.RdData_98(out_reg_r_98),
.RdData_99(out_reg_r_99),
.RdData_100(out_reg_r_100),
.RdData_101(out_reg_r_101),
.RdData_102(out_reg_r_102),
.RdData_103(out_reg_r_103),
.RdData_104(out_reg_r_104),
.RdData_105(out_reg_r_105),
.RdData_106(out_reg_r_106),
.RdData_107(out_reg_r_107),
.RdData_108(out_reg_r_108),
.RdData_109(out_reg_r_109),
.RdData_110(out_reg_r_110),
.RdData_111(out_reg_r_111),
.RdData_112(out_reg_r_112),
.RdData_113(out_reg_r_113),
.RdData_114(out_reg_r_114),
.RdData_115(out_reg_r_115),
.RdData_116(out_reg_r_116),
.RdData_117(out_reg_r_117),
.RdData_118(out_reg_r_118),
.RdData_119(out_reg_r_119),
.RdData_120(out_reg_r_120),
.RdData_121(out_reg_r_121),
.RdData_122(out_reg_r_122),
.RdData_123(out_reg_r_123),
.RdData_124(out_reg_r_124),
.RdData_125(out_reg_r_125),
.RdData_126(out_reg_r_126),
.RdData_127(out_reg_r_127)

);





Reg_File #(.BITS(BITS),.NUMBER_OF_REGISTERS(NUMBER_OF_ENABLE_BITS)) Reg_File_IMG 
( 

.WrEn(reg_en) , 
.clk(clk) ,
.rst(rst) , 
  
.WrData_0(memory_imag_output_0),
.WrData_1(memory_imag_output_0),
.WrData_2(memory_imag_output_0),
.WrData_3(memory_imag_output_0),
.WrData_4(memory_imag_output_1),
.WrData_5(memory_imag_output_1),
.WrData_6(memory_imag_output_1),
.WrData_7(memory_imag_output_1),
.WrData_8(memory_imag_output_2),
.WrData_9(memory_imag_output_2),
.WrData_10(memory_imag_output_2),
.WrData_11(memory_imag_output_2),
.WrData_12(memory_imag_output_3),
.WrData_13(memory_imag_output_3),
.WrData_14(memory_imag_output_3),
.WrData_15(memory_imag_output_3),
.WrData_16(memory_imag_output_4),
.WrData_17(memory_imag_output_4),
.WrData_18(memory_imag_output_4),
.WrData_19(memory_imag_output_4),
.WrData_20(memory_imag_output_5),
.WrData_21(memory_imag_output_5),
.WrData_22(memory_imag_output_5),
.WrData_23(memory_imag_output_5),
.WrData_24(memory_imag_output_6),
.WrData_25(memory_imag_output_6),
.WrData_26(memory_imag_output_6),
.WrData_27(memory_imag_output_6),
.WrData_28(memory_imag_output_7),
.WrData_29(memory_imag_output_7),
.WrData_30(memory_imag_output_7),
.WrData_31(memory_imag_output_7),
.WrData_32(memory_imag_output_8),
.WrData_33(memory_imag_output_8),
.WrData_34(memory_imag_output_8),
.WrData_35(memory_imag_output_8),
.WrData_36(memory_imag_output_9),
.WrData_37(memory_imag_output_9),
.WrData_38(memory_imag_output_9),
.WrData_39(memory_imag_output_9),
.WrData_40(memory_imag_output_10),
.WrData_41(memory_imag_output_10),
.WrData_42(memory_imag_output_10),
.WrData_43(memory_imag_output_10),
.WrData_44(memory_imag_output_11),
.WrData_45(memory_imag_output_11),
.WrData_46(memory_imag_output_11),
.WrData_47(memory_imag_output_11),
.WrData_48(memory_imag_output_12),
.WrData_49(memory_imag_output_12),
.WrData_50(memory_imag_output_12),
.WrData_51(memory_imag_output_12),
.WrData_52(memory_imag_output_13),
.WrData_53(memory_imag_output_13),
.WrData_54(memory_imag_output_13),
.WrData_55(memory_imag_output_13),
.WrData_56(memory_imag_output_14),
.WrData_57(memory_imag_output_14),
.WrData_58(memory_imag_output_14),
.WrData_59(memory_imag_output_14),
.WrData_60(memory_imag_output_15),
.WrData_61(memory_imag_output_15),
.WrData_62(memory_imag_output_15),
.WrData_63(memory_imag_output_15),
.WrData_64(memory_imag_output_16),
.WrData_65(memory_imag_output_16),
.WrData_66(memory_imag_output_16),
.WrData_67(memory_imag_output_16),
.WrData_68(memory_imag_output_17),
.WrData_69(memory_imag_output_17),
.WrData_70(memory_imag_output_17),
.WrData_71(memory_imag_output_17),
.WrData_72(memory_imag_output_18),
.WrData_73(memory_imag_output_18),
.WrData_74(memory_imag_output_18),
.WrData_75(memory_imag_output_18),
.WrData_76(memory_imag_output_19),
.WrData_77(memory_imag_output_19),
.WrData_78(memory_imag_output_19),
.WrData_79(memory_imag_output_19),
.WrData_80(memory_imag_output_20),
.WrData_81(memory_imag_output_20),
.WrData_82(memory_imag_output_20),
.WrData_83(memory_imag_output_20),
.WrData_84(memory_imag_output_21),
.WrData_85(memory_imag_output_21),
.WrData_86(memory_imag_output_21),
.WrData_87(memory_imag_output_21),
.WrData_88(memory_imag_output_22),
.WrData_89(memory_imag_output_22),
.WrData_90(memory_imag_output_22),
.WrData_91(memory_imag_output_22),
.WrData_92(memory_imag_output_23),
.WrData_93(memory_imag_output_23),
.WrData_94(memory_imag_output_23),
.WrData_95(memory_imag_output_23),
.WrData_96(memory_imag_output_24),
.WrData_97(memory_imag_output_24),
.WrData_98(memory_imag_output_24),
.WrData_99(memory_imag_output_24),
.WrData_100(memory_imag_output_25),
.WrData_101(memory_imag_output_25),
.WrData_102(memory_imag_output_25),
.WrData_103(memory_imag_output_25),
.WrData_104(memory_imag_output_26),
.WrData_105(memory_imag_output_26),
.WrData_106(memory_imag_output_26),
.WrData_107(memory_imag_output_26),
.WrData_108(memory_imag_output_27),
.WrData_109(memory_imag_output_27),
.WrData_110(memory_imag_output_27),
.WrData_111(memory_imag_output_27),
.WrData_112(memory_imag_output_28),
.WrData_113(memory_imag_output_28),
.WrData_114(memory_imag_output_28),
.WrData_115(memory_imag_output_28),
.WrData_116(memory_imag_output_29),
.WrData_117(memory_imag_output_29),
.WrData_118(memory_imag_output_29),
.WrData_119(memory_imag_output_29),
.WrData_120(memory_imag_output_30),
.WrData_121(memory_imag_output_30),
.WrData_122(memory_imag_output_30),
.WrData_123(memory_imag_output_30),
.WrData_124(memory_imag_output_31),
.WrData_125(memory_imag_output_31),
.WrData_126(memory_imag_output_31),
.WrData_127(memory_imag_output_31),


.RdData_0(out_reg_i_0),
.RdData_1(out_reg_i_1),
.RdData_2(out_reg_i_2),
.RdData_3(out_reg_i_3),
.RdData_4(out_reg_i_4),
.RdData_5(out_reg_i_5),
.RdData_6(out_reg_i_6),
.RdData_7(out_reg_i_7),
.RdData_8(out_reg_i_8),
.RdData_9(out_reg_i_9),
.RdData_10(out_reg_i_10),
.RdData_11(out_reg_i_11),
.RdData_12(out_reg_i_12),
.RdData_13(out_reg_i_13),
.RdData_14(out_reg_i_14),
.RdData_15(out_reg_i_15),
.RdData_16(out_reg_i_16),
.RdData_17(out_reg_i_17),
.RdData_18(out_reg_i_18),
.RdData_19(out_reg_i_19),
.RdData_20(out_reg_i_20),
.RdData_21(out_reg_i_21),
.RdData_22(out_reg_i_22),
.RdData_23(out_reg_i_23),
.RdData_24(out_reg_i_24),
.RdData_25(out_reg_i_25),
.RdData_26(out_reg_i_26),
.RdData_27(out_reg_i_27),
.RdData_28(out_reg_i_28),
.RdData_29(out_reg_i_29),
.RdData_30(out_reg_i_30),
.RdData_31(out_reg_i_31),
.RdData_32(out_reg_i_32),
.RdData_33(out_reg_i_33),
.RdData_34(out_reg_i_34),
.RdData_35(out_reg_i_35),
.RdData_36(out_reg_i_36),
.RdData_37(out_reg_i_37),
.RdData_38(out_reg_i_38),
.RdData_39(out_reg_i_39),
.RdData_40(out_reg_i_40),
.RdData_41(out_reg_i_41),
.RdData_42(out_reg_i_42),
.RdData_43(out_reg_i_43),
.RdData_44(out_reg_i_44),
.RdData_45(out_reg_i_45),
.RdData_46(out_reg_i_46),
.RdData_47(out_reg_i_47),
.RdData_48(out_reg_i_48),
.RdData_49(out_reg_i_49),
.RdData_50(out_reg_i_50),
.RdData_51(out_reg_i_51),
.RdData_52(out_reg_i_52),
.RdData_53(out_reg_i_53),
.RdData_54(out_reg_i_54),
.RdData_55(out_reg_i_55),
.RdData_56(out_reg_i_56),
.RdData_57(out_reg_i_57),
.RdData_58(out_reg_i_58),
.RdData_59(out_reg_i_59),
.RdData_60(out_reg_i_60),
.RdData_61(out_reg_i_61),
.RdData_62(out_reg_i_62),
.RdData_63(out_reg_i_63),
.RdData_64(out_reg_i_64),
.RdData_65(out_reg_i_65),
.RdData_66(out_reg_i_66),
.RdData_67(out_reg_i_67),
.RdData_68(out_reg_i_68),
.RdData_69(out_reg_i_69),
.RdData_70(out_reg_i_70),
.RdData_71(out_reg_i_71),
.RdData_72(out_reg_i_72),
.RdData_73(out_reg_i_73),
.RdData_74(out_reg_i_74),
.RdData_75(out_reg_i_75),
.RdData_76(out_reg_i_76),
.RdData_77(out_reg_i_77),
.RdData_78(out_reg_i_78),
.RdData_79(out_reg_i_79),
.RdData_80(out_reg_i_80),
.RdData_81(out_reg_i_81),
.RdData_82(out_reg_i_82),
.RdData_83(out_reg_i_83),
.RdData_84(out_reg_i_84),
.RdData_85(out_reg_i_85),
.RdData_86(out_reg_i_86),
.RdData_87(out_reg_i_87),
.RdData_88(out_reg_i_88),
.RdData_89(out_reg_i_89),
.RdData_90(out_reg_i_90),
.RdData_91(out_reg_i_91),
.RdData_92(out_reg_i_92),
.RdData_93(out_reg_i_93),
.RdData_94(out_reg_i_94),
.RdData_95(out_reg_i_95),
.RdData_96(out_reg_i_96),
.RdData_97(out_reg_i_97),
.RdData_98(out_reg_i_98),
.RdData_99(out_reg_i_99),
.RdData_100(out_reg_i_100),
.RdData_101(out_reg_i_101),
.RdData_102(out_reg_i_102),
.RdData_103(out_reg_i_103),
.RdData_104(out_reg_i_104),
.RdData_105(out_reg_i_105),
.RdData_106(out_reg_i_106),
.RdData_107(out_reg_i_107),
.RdData_108(out_reg_i_108),
.RdData_109(out_reg_i_109),
.RdData_110(out_reg_i_110),
.RdData_111(out_reg_i_111),
.RdData_112(out_reg_i_112),
.RdData_113(out_reg_i_113),
.RdData_114(out_reg_i_114),
.RdData_115(out_reg_i_115),
.RdData_116(out_reg_i_116),
.RdData_117(out_reg_i_117),
.RdData_118(out_reg_i_118),
.RdData_119(out_reg_i_119),
.RdData_120(out_reg_i_120),
.RdData_121(out_reg_i_121),
.RdData_122(out_reg_i_122),
.RdData_123(out_reg_i_123),
.RdData_124(out_reg_i_124),
.RdData_125(out_reg_i_125),
.RdData_126(out_reg_i_126),
.RdData_127(out_reg_i_127)

);





Reg_File_64 #(.BITS(BITS),.NUMBER_OF_REGISTERS(64)) Reg_File_twiddle_real
(
.WrEn(twiddle_reg_en) , 
.clk(clk) ,
.rst(rst) , 

.WrData_0(ROM_out_twiddle_r_0),
.WrData_1(ROM_out_twiddle_r_0),
.WrData_2(ROM_out_twiddle_r_0),
.WrData_3(ROM_out_twiddle_r_0),
.WrData_4(ROM_out_twiddle_r_1),
.WrData_5(ROM_out_twiddle_r_1),
.WrData_6(ROM_out_twiddle_r_1),
.WrData_7(ROM_out_twiddle_r_1),
.WrData_8(ROM_out_twiddle_r_2),
.WrData_9(ROM_out_twiddle_r_2),
.WrData_10(ROM_out_twiddle_r_2),
.WrData_11(ROM_out_twiddle_r_2),
.WrData_12(ROM_out_twiddle_r_3),
.WrData_13(ROM_out_twiddle_r_3),
.WrData_14(ROM_out_twiddle_r_3),
.WrData_15(ROM_out_twiddle_r_3),
.WrData_16(ROM_out_twiddle_r_4),
.WrData_17(ROM_out_twiddle_r_4),
.WrData_18(ROM_out_twiddle_r_4),
.WrData_19(ROM_out_twiddle_r_4),
.WrData_20(ROM_out_twiddle_r_5),
.WrData_21(ROM_out_twiddle_r_5),
.WrData_22(ROM_out_twiddle_r_5),
.WrData_23(ROM_out_twiddle_r_5),
.WrData_24(ROM_out_twiddle_r_6),
.WrData_25(ROM_out_twiddle_r_6),
.WrData_26(ROM_out_twiddle_r_6),
.WrData_27(ROM_out_twiddle_r_6),
.WrData_28(ROM_out_twiddle_r_7),
.WrData_29(ROM_out_twiddle_r_7),
.WrData_30(ROM_out_twiddle_r_7),
.WrData_31(ROM_out_twiddle_r_7),
.WrData_32(ROM_out_twiddle_r_8),
.WrData_33(ROM_out_twiddle_r_8),
.WrData_34(ROM_out_twiddle_r_8),
.WrData_35(ROM_out_twiddle_r_8),
.WrData_36(ROM_out_twiddle_r_9),
.WrData_37(ROM_out_twiddle_r_9),
.WrData_38(ROM_out_twiddle_r_9),
.WrData_39(ROM_out_twiddle_r_9),
.WrData_40(ROM_out_twiddle_r_10),
.WrData_41(ROM_out_twiddle_r_10),
.WrData_42(ROM_out_twiddle_r_10),
.WrData_43(ROM_out_twiddle_r_10),
.WrData_44(ROM_out_twiddle_r_11),
.WrData_45(ROM_out_twiddle_r_11),
.WrData_46(ROM_out_twiddle_r_11),
.WrData_47(ROM_out_twiddle_r_11),
.WrData_48(ROM_out_twiddle_r_12),
.WrData_49(ROM_out_twiddle_r_12),
.WrData_50(ROM_out_twiddle_r_12),
.WrData_51(ROM_out_twiddle_r_12),
.WrData_52(ROM_out_twiddle_r_13),
.WrData_53(ROM_out_twiddle_r_13),
.WrData_54(ROM_out_twiddle_r_13),
.WrData_55(ROM_out_twiddle_r_13),
.WrData_56(ROM_out_twiddle_r_14),
.WrData_57(ROM_out_twiddle_r_14),
.WrData_58(ROM_out_twiddle_r_14),
.WrData_59(ROM_out_twiddle_r_14),
.WrData_60(ROM_out_twiddle_r_15),
.WrData_61(ROM_out_twiddle_r_15),
.WrData_62(ROM_out_twiddle_r_15),
.WrData_63(ROM_out_twiddle_r_15),


.RdData_0(out_reg_twiddle_r_0),
.RdData_1(out_reg_twiddle_r_1),
.RdData_2(out_reg_twiddle_r_2),
.RdData_3(out_reg_twiddle_r_3),
.RdData_4(out_reg_twiddle_r_4),
.RdData_5(out_reg_twiddle_r_5),
.RdData_6(out_reg_twiddle_r_6),
.RdData_7(out_reg_twiddle_r_7),
.RdData_8(out_reg_twiddle_r_8),
.RdData_9(out_reg_twiddle_r_9),
.RdData_10(out_reg_twiddle_r_10),
.RdData_11(out_reg_twiddle_r_11),
.RdData_12(out_reg_twiddle_r_12),
.RdData_13(out_reg_twiddle_r_13),
.RdData_14(out_reg_twiddle_r_14),
.RdData_15(out_reg_twiddle_r_15),
.RdData_16(out_reg_twiddle_r_16),
.RdData_17(out_reg_twiddle_r_17),
.RdData_18(out_reg_twiddle_r_18),
.RdData_19(out_reg_twiddle_r_19),
.RdData_20(out_reg_twiddle_r_20),
.RdData_21(out_reg_twiddle_r_21),
.RdData_22(out_reg_twiddle_r_22),
.RdData_23(out_reg_twiddle_r_23),
.RdData_24(out_reg_twiddle_r_24),
.RdData_25(out_reg_twiddle_r_25),
.RdData_26(out_reg_twiddle_r_26),
.RdData_27(out_reg_twiddle_r_27),
.RdData_28(out_reg_twiddle_r_28),
.RdData_29(out_reg_twiddle_r_29),
.RdData_30(out_reg_twiddle_r_30),
.RdData_31(out_reg_twiddle_r_31),
.RdData_32(out_reg_twiddle_r_32),
.RdData_33(out_reg_twiddle_r_33),
.RdData_34(out_reg_twiddle_r_34),
.RdData_35(out_reg_twiddle_r_35),
.RdData_36(out_reg_twiddle_r_36),
.RdData_37(out_reg_twiddle_r_37),
.RdData_38(out_reg_twiddle_r_38),
.RdData_39(out_reg_twiddle_r_39),
.RdData_40(out_reg_twiddle_r_40),
.RdData_41(out_reg_twiddle_r_41),
.RdData_42(out_reg_twiddle_r_42),
.RdData_43(out_reg_twiddle_r_43),
.RdData_44(out_reg_twiddle_r_44),
.RdData_45(out_reg_twiddle_r_45),
.RdData_46(out_reg_twiddle_r_46),
.RdData_47(out_reg_twiddle_r_47),
.RdData_48(out_reg_twiddle_r_48),
.RdData_49(out_reg_twiddle_r_49),
.RdData_50(out_reg_twiddle_r_50),
.RdData_51(out_reg_twiddle_r_51),
.RdData_52(out_reg_twiddle_r_52),
.RdData_53(out_reg_twiddle_r_53),
.RdData_54(out_reg_twiddle_r_54),
.RdData_55(out_reg_twiddle_r_55),
.RdData_56(out_reg_twiddle_r_56),
.RdData_57(out_reg_twiddle_r_57),
.RdData_58(out_reg_twiddle_r_58),
.RdData_59(out_reg_twiddle_r_59),
.RdData_60(out_reg_twiddle_r_60),
.RdData_61(out_reg_twiddle_r_61),
.RdData_62(out_reg_twiddle_r_62),
.RdData_63(out_reg_twiddle_r_63)

);








Reg_File_64 #(.BITS(BITS),.NUMBER_OF_REGISTERS(64)) Reg_File_twiddle_img
(
.WrEn(twiddle_reg_en) , 
.clk(clk) ,
.rst(rst) , 

.WrData_0(ROM_out_twiddle_i_0),
.WrData_1(ROM_out_twiddle_i_0),
.WrData_2(ROM_out_twiddle_i_0),
.WrData_3(ROM_out_twiddle_i_0),
.WrData_4(ROM_out_twiddle_i_1),
.WrData_5(ROM_out_twiddle_i_1),
.WrData_6(ROM_out_twiddle_i_1),
.WrData_7(ROM_out_twiddle_i_1),
.WrData_8(ROM_out_twiddle_i_2),
.WrData_9(ROM_out_twiddle_i_2),
.WrData_10(ROM_out_twiddle_i_2),
.WrData_11(ROM_out_twiddle_i_2),
.WrData_12(ROM_out_twiddle_i_3),
.WrData_13(ROM_out_twiddle_i_3),
.WrData_14(ROM_out_twiddle_i_3),
.WrData_15(ROM_out_twiddle_i_3),
.WrData_16(ROM_out_twiddle_i_4),
.WrData_17(ROM_out_twiddle_i_4),
.WrData_18(ROM_out_twiddle_i_4),
.WrData_19(ROM_out_twiddle_i_4),
.WrData_20(ROM_out_twiddle_i_5),
.WrData_21(ROM_out_twiddle_i_5),
.WrData_22(ROM_out_twiddle_i_5),
.WrData_23(ROM_out_twiddle_i_5),
.WrData_24(ROM_out_twiddle_i_6),
.WrData_25(ROM_out_twiddle_i_6),
.WrData_26(ROM_out_twiddle_i_6),
.WrData_27(ROM_out_twiddle_i_6),
.WrData_28(ROM_out_twiddle_i_7),
.WrData_29(ROM_out_twiddle_i_7),
.WrData_30(ROM_out_twiddle_i_7),
.WrData_31(ROM_out_twiddle_i_7),
.WrData_32(ROM_out_twiddle_i_8),
.WrData_33(ROM_out_twiddle_i_8),
.WrData_34(ROM_out_twiddle_i_8),
.WrData_35(ROM_out_twiddle_i_8),
.WrData_36(ROM_out_twiddle_i_9),
.WrData_37(ROM_out_twiddle_i_9),
.WrData_38(ROM_out_twiddle_i_9),
.WrData_39(ROM_out_twiddle_i_9),
.WrData_40(ROM_out_twiddle_i_10),
.WrData_41(ROM_out_twiddle_i_10),
.WrData_42(ROM_out_twiddle_i_10),
.WrData_43(ROM_out_twiddle_i_10),
.WrData_44(ROM_out_twiddle_i_11),
.WrData_45(ROM_out_twiddle_i_11),
.WrData_46(ROM_out_twiddle_i_11),
.WrData_47(ROM_out_twiddle_i_11),
.WrData_48(ROM_out_twiddle_i_12),
.WrData_49(ROM_out_twiddle_i_12),
.WrData_50(ROM_out_twiddle_i_12),
.WrData_51(ROM_out_twiddle_i_12),
.WrData_52(ROM_out_twiddle_i_13),
.WrData_53(ROM_out_twiddle_i_13),
.WrData_54(ROM_out_twiddle_i_13),
.WrData_55(ROM_out_twiddle_i_13),
.WrData_56(ROM_out_twiddle_i_14),
.WrData_57(ROM_out_twiddle_i_14),
.WrData_58(ROM_out_twiddle_i_14),
.WrData_59(ROM_out_twiddle_i_14),
.WrData_60(ROM_out_twiddle_i_15),
.WrData_61(ROM_out_twiddle_i_15),
.WrData_62(ROM_out_twiddle_i_15),
.WrData_63(ROM_out_twiddle_i_15),


.RdData_0(out_reg_twiddle_i_0),
.RdData_1(out_reg_twiddle_i_1),
.RdData_2(out_reg_twiddle_i_2),
.RdData_3(out_reg_twiddle_i_3),
.RdData_4(out_reg_twiddle_i_4),
.RdData_5(out_reg_twiddle_i_5),
.RdData_6(out_reg_twiddle_i_6),
.RdData_7(out_reg_twiddle_i_7),
.RdData_8(out_reg_twiddle_i_8),
.RdData_9(out_reg_twiddle_i_9),
.RdData_10(out_reg_twiddle_i_10),
.RdData_11(out_reg_twiddle_i_11),
.RdData_12(out_reg_twiddle_i_12),
.RdData_13(out_reg_twiddle_i_13),
.RdData_14(out_reg_twiddle_i_14),
.RdData_15(out_reg_twiddle_i_15),
.RdData_16(out_reg_twiddle_i_16),
.RdData_17(out_reg_twiddle_i_17),
.RdData_18(out_reg_twiddle_i_18),
.RdData_19(out_reg_twiddle_i_19),
.RdData_20(out_reg_twiddle_i_20),
.RdData_21(out_reg_twiddle_i_21),
.RdData_22(out_reg_twiddle_i_22),
.RdData_23(out_reg_twiddle_i_23),
.RdData_24(out_reg_twiddle_i_24),
.RdData_25(out_reg_twiddle_i_25),
.RdData_26(out_reg_twiddle_i_26),
.RdData_27(out_reg_twiddle_i_27),
.RdData_28(out_reg_twiddle_i_28),
.RdData_29(out_reg_twiddle_i_29),
.RdData_30(out_reg_twiddle_i_30),
.RdData_31(out_reg_twiddle_i_31),
.RdData_32(out_reg_twiddle_i_32),
.RdData_33(out_reg_twiddle_i_33),
.RdData_34(out_reg_twiddle_i_34),
.RdData_35(out_reg_twiddle_i_35),
.RdData_36(out_reg_twiddle_i_36),
.RdData_37(out_reg_twiddle_i_37),
.RdData_38(out_reg_twiddle_i_38),
.RdData_39(out_reg_twiddle_i_39),
.RdData_40(out_reg_twiddle_i_40),
.RdData_41(out_reg_twiddle_i_41),
.RdData_42(out_reg_twiddle_i_42),
.RdData_43(out_reg_twiddle_i_43),
.RdData_44(out_reg_twiddle_i_44),
.RdData_45(out_reg_twiddle_i_45),
.RdData_46(out_reg_twiddle_i_46),
.RdData_47(out_reg_twiddle_i_47),
.RdData_48(out_reg_twiddle_i_48),
.RdData_49(out_reg_twiddle_i_49),
.RdData_50(out_reg_twiddle_i_50),
.RdData_51(out_reg_twiddle_i_51),
.RdData_52(out_reg_twiddle_i_52),
.RdData_53(out_reg_twiddle_i_53),
.RdData_54(out_reg_twiddle_i_54),
.RdData_55(out_reg_twiddle_i_55),
.RdData_56(out_reg_twiddle_i_56),
.RdData_57(out_reg_twiddle_i_57),
.RdData_58(out_reg_twiddle_i_58),
.RdData_59(out_reg_twiddle_i_59),
.RdData_60(out_reg_twiddle_i_60),
.RdData_61(out_reg_twiddle_i_61),
.RdData_62(out_reg_twiddle_i_62),
.RdData_63(out_reg_twiddle_i_63)

);









Butterfly_Column_Top #(.BITS(BITS)) unt
(
.rst(rst),
//.clk(clk_4),
.t0_r(out_reg_r_0),
.t1_r(out_reg_r_1),
.t2_r(out_reg_r_2),
.t3_r(out_reg_r_3),
.t4_r(out_reg_r_4),
.t5_r(out_reg_r_5),
.t6_r(out_reg_r_6),
.t7_r(out_reg_r_7),
.t8_r(out_reg_r_8),
.t9_r(out_reg_r_9),
.t10_r(out_reg_r_10),
.t11_r(out_reg_r_11),
.t12_r(out_reg_r_12),
.t13_r(out_reg_r_13),
.t14_r(out_reg_r_14),
.t15_r(out_reg_r_15),
.t16_r(out_reg_r_16),
.t17_r(out_reg_r_17),
.t18_r(out_reg_r_18),
.t19_r(out_reg_r_19),
.t20_r(out_reg_r_20),
.t21_r(out_reg_r_21),
.t22_r(out_reg_r_22),
.t23_r(out_reg_r_23),
.t24_r(out_reg_r_24),
.t25_r(out_reg_r_25),
.t26_r(out_reg_r_26),
.t27_r(out_reg_r_27),
.t28_r(out_reg_r_28),
.t29_r(out_reg_r_29),
.t30_r(out_reg_r_30),
.t31_r(out_reg_r_31),
.t32_r(out_reg_r_32),
.t33_r(out_reg_r_33),
.t34_r(out_reg_r_34),
.t35_r(out_reg_r_35),
.t36_r(out_reg_r_36),
.t37_r(out_reg_r_37),
.t38_r(out_reg_r_38),
.t39_r(out_reg_r_39),
.t40_r(out_reg_r_40),
.t41_r(out_reg_r_41),
.t42_r(out_reg_r_42),
.t43_r(out_reg_r_43),
.t44_r(out_reg_r_44),
.t45_r(out_reg_r_45),
.t46_r(out_reg_r_46),
.t47_r(out_reg_r_47),
.t48_r(out_reg_r_48),
.t49_r(out_reg_r_49),
.t50_r(out_reg_r_50),
.t51_r(out_reg_r_51),
.t52_r(out_reg_r_52),
.t53_r(out_reg_r_53),
.t54_r(out_reg_r_54),
.t55_r(out_reg_r_55),
.t56_r(out_reg_r_56),
.t57_r(out_reg_r_57),
.t58_r(out_reg_r_58),
.t59_r(out_reg_r_59),
.t60_r(out_reg_r_60),
.t61_r(out_reg_r_61),
.t62_r(out_reg_r_62),
.t63_r(out_reg_r_63),
.t64_r(out_reg_r_64),
.t65_r(out_reg_r_65),
.t66_r(out_reg_r_66),
.t67_r(out_reg_r_67),
.t68_r(out_reg_r_68),
.t69_r(out_reg_r_69),
.t70_r(out_reg_r_70),
.t71_r(out_reg_r_71),
.t72_r(out_reg_r_72),
.t73_r(out_reg_r_73),
.t74_r(out_reg_r_74),
.t75_r(out_reg_r_75),
.t76_r(out_reg_r_76),
.t77_r(out_reg_r_77),
.t78_r(out_reg_r_78),
.t79_r(out_reg_r_79),
.t80_r(out_reg_r_80),
.t81_r(out_reg_r_81),
.t82_r(out_reg_r_82),
.t83_r(out_reg_r_83),
.t84_r(out_reg_r_84),
.t85_r(out_reg_r_85),
.t86_r(out_reg_r_86),
.t87_r(out_reg_r_87),
.t88_r(out_reg_r_88),
.t89_r(out_reg_r_89),
.t90_r(out_reg_r_90),
.t91_r(out_reg_r_91),
.t92_r(out_reg_r_92),
.t93_r(out_reg_r_93),
.t94_r(out_reg_r_94),
.t95_r(out_reg_r_95),
.t96_r(out_reg_r_96),
.t97_r(out_reg_r_97),
.t98_r(out_reg_r_98),
.t99_r(out_reg_r_99),
.t100_r(out_reg_r_100),
.t101_r(out_reg_r_101),
.t102_r(out_reg_r_102),
.t103_r(out_reg_r_103),
.t104_r(out_reg_r_104),
.t105_r(out_reg_r_105),
.t106_r(out_reg_r_106),
.t107_r(out_reg_r_107),
.t108_r(out_reg_r_108),
.t109_r(out_reg_r_109),
.t110_r(out_reg_r_110),
.t111_r(out_reg_r_111),
.t112_r(out_reg_r_112),
.t113_r(out_reg_r_113),
.t114_r(out_reg_r_114),
.t115_r(out_reg_r_115),
.t116_r(out_reg_r_116),
.t117_r(out_reg_r_117),
.t118_r(out_reg_r_118),
.t119_r(out_reg_r_119),
.t120_r(out_reg_r_120),
.t121_r(out_reg_r_121),
.t122_r(out_reg_r_122),
.t123_r(out_reg_r_123),
.t124_r(out_reg_r_124),
.t125_r(out_reg_r_125),
.t126_r(out_reg_r_126),
.t127_r(out_reg_r_127),


.t0_i(out_reg_i_0),
.t1_i(out_reg_i_1),
.t2_i(out_reg_i_2),
.t3_i(out_reg_i_3),
.t4_i(out_reg_i_4),
.t5_i(out_reg_i_5),
.t6_i(out_reg_i_6),
.t7_i(out_reg_i_7),
.t8_i(out_reg_i_8),
.t9_i(out_reg_i_9),
.t10_i(out_reg_i_10),
.t11_i(out_reg_i_11),
.t12_i(out_reg_i_12),
.t13_i(out_reg_i_13),
.t14_i(out_reg_i_14),
.t15_i(out_reg_i_15),
.t16_i(out_reg_i_16),
.t17_i(out_reg_i_17),
.t18_i(out_reg_i_18),
.t19_i(out_reg_i_19),
.t20_i(out_reg_i_20),
.t21_i(out_reg_i_21),
.t22_i(out_reg_i_22),
.t23_i(out_reg_i_23),
.t24_i(out_reg_i_24),
.t25_i(out_reg_i_25),
.t26_i(out_reg_i_26),
.t27_i(out_reg_i_27),
.t28_i(out_reg_i_28),
.t29_i(out_reg_i_29),
.t30_i(out_reg_i_30),
.t31_i(out_reg_i_31),
.t32_i(out_reg_i_32),
.t33_i(out_reg_i_33),
.t34_i(out_reg_i_34),
.t35_i(out_reg_i_35),
.t36_i(out_reg_i_36),
.t37_i(out_reg_i_37),
.t38_i(out_reg_i_38),
.t39_i(out_reg_i_39),
.t40_i(out_reg_i_40),
.t41_i(out_reg_i_41),
.t42_i(out_reg_i_42),
.t43_i(out_reg_i_43),
.t44_i(out_reg_i_44),
.t45_i(out_reg_i_45),
.t46_i(out_reg_i_46),
.t47_i(out_reg_i_47),
.t48_i(out_reg_i_48),
.t49_i(out_reg_i_49),
.t50_i(out_reg_i_50),
.t51_i(out_reg_i_51),
.t52_i(out_reg_i_52),
.t53_i(out_reg_i_53),
.t54_i(out_reg_i_54),
.t55_i(out_reg_i_55),
.t56_i(out_reg_i_56),
.t57_i(out_reg_i_57),
.t58_i(out_reg_i_58),
.t59_i(out_reg_i_59),
.t60_i(out_reg_i_60),
.t61_i(out_reg_i_61),
.t62_i(out_reg_i_62),
.t63_i(out_reg_i_63),
.t64_i(out_reg_i_64),
.t65_i(out_reg_i_65),
.t66_i(out_reg_i_66),
.t67_i(out_reg_i_67),
.t68_i(out_reg_i_68),
.t69_i(out_reg_i_69),
.t70_i(out_reg_i_70),
.t71_i(out_reg_i_71),
.t72_i(out_reg_i_72),
.t73_i(out_reg_i_73),
.t74_i(out_reg_i_74),
.t75_i(out_reg_i_75),
.t76_i(out_reg_i_76),
.t77_i(out_reg_i_77),
.t78_i(out_reg_i_78),
.t79_i(out_reg_i_79),
.t80_i(out_reg_i_80),
.t81_i(out_reg_i_81),
.t82_i(out_reg_i_82),
.t83_i(out_reg_i_83),
.t84_i(out_reg_i_84),
.t85_i(out_reg_i_85),
.t86_i(out_reg_i_86),
.t87_i(out_reg_i_87),
.t88_i(out_reg_i_88),
.t89_i(out_reg_i_89),
.t90_i(out_reg_i_90),
.t91_i(out_reg_i_91),
.t92_i(out_reg_i_92),
.t93_i(out_reg_i_93),
.t94_i(out_reg_i_94),
.t95_i(out_reg_i_95),
.t96_i(out_reg_i_96),
.t97_i(out_reg_i_97),
.t98_i(out_reg_i_98),
.t99_i(out_reg_i_99),
.t100_i(out_reg_i_100),
.t101_i(out_reg_i_101),
.t102_i(out_reg_i_102),
.t103_i(out_reg_i_103),
.t104_i(out_reg_i_104),
.t105_i(out_reg_i_105),
.t106_i(out_reg_i_106),
.t107_i(out_reg_i_107),
.t108_i(out_reg_i_108),
.t109_i(out_reg_i_109),
.t110_i(out_reg_i_110),
.t111_i(out_reg_i_111),
.t112_i(out_reg_i_112),
.t113_i(out_reg_i_113),
.t114_i(out_reg_i_114),
.t115_i(out_reg_i_115),
.t116_i(out_reg_i_116),
.t117_i(out_reg_i_117),
.t118_i(out_reg_i_118),
.t119_i(out_reg_i_119),
.t120_i(out_reg_i_120),
.t121_i(out_reg_i_121),
.t122_i(out_reg_i_122),
.t123_i(out_reg_i_123),
.t124_i(out_reg_i_124),
.t125_i(out_reg_i_125),
.t126_i(out_reg_i_126),
.t127_i(out_reg_i_127),




.s0_r(s0_r),
.s0_i(s0_i),
.s1_r(s1_r),
.s1_i(s1_i),
.s2_r(s2_r),
.s2_i(s2_i),
.s3_r(s3_r),
.s3_i(s3_i),
.s4_r(s4_r),
.s4_i(s4_i),
.s5_r(s5_r),
.s5_i(s5_i),
.s6_r(s6_r),
.s6_i(s6_i),
.s7_r(s7_r),
.s7_i(s7_i),
.s8_r(s8_r),
.s8_i(s8_i),
.s9_r(s9_r),
.s9_i(s9_i),
.s10_r(s10_r),
.s10_i(s10_i),
.s11_r(s11_r),
.s11_i(s11_i),
.s12_r(s12_r),
.s12_i(s12_i),
.s13_r(s13_r),
.s13_i(s13_i),
.s14_r(s14_r),
.s14_i(s14_i),
.s15_r(s15_r),
.s15_i(s15_i),
.s16_r(s16_r),
.s16_i(s16_i),
.s17_r(s17_r),
.s17_i(s17_i),
.s18_r(s18_r),
.s18_i(s18_i),
.s19_r(s19_r),
.s19_i(s19_i),
.s20_r(s20_r),
.s20_i(s20_i),
.s21_r(s21_r),
.s21_i(s21_i),
.s22_r(s22_r),
.s22_i(s22_i),
.s23_r(s23_r),
.s23_i(s23_i),
.s24_r(s24_r),
.s24_i(s24_i),
.s25_r(s25_r),
.s25_i(s25_i),
.s26_r(s26_r),
.s26_i(s26_i),
.s27_r(s27_r),
.s27_i(s27_i),
.s28_r(s28_r),
.s28_i(s28_i),
.s29_r(s29_r),
.s29_i(s29_i),
.s30_r(s30_r),
.s30_i(s30_i),
.s31_r(s31_r),
.s31_i(s31_i),
.s32_r(s32_r),
.s32_i(s32_i),
.s33_r(s33_r),
.s33_i(s33_i),
.s34_r(s34_r),
.s34_i(s34_i),
.s35_r(s35_r),
.s35_i(s35_i),
.s36_r(s36_r),
.s36_i(s36_i),
.s37_r(s37_r),
.s37_i(s37_i),
.s38_r(s38_r),
.s38_i(s38_i),
.s39_r(s39_r),
.s39_i(s39_i),
.s40_r(s40_r),
.s40_i(s40_i),
.s41_r(s41_r),
.s41_i(s41_i),
.s42_r(s42_r),
.s42_i(s42_i),
.s43_r(s43_r),
.s43_i(s43_i),
.s44_r(s44_r),
.s44_i(s44_i),
.s45_r(s45_r),
.s45_i(s45_i),
.s46_r(s46_r),
.s46_i(s46_i),
.s47_r(s47_r),
.s47_i(s47_i),
.s48_r(s48_r),
.s48_i(s48_i),
.s49_r(s49_r),
.s49_i(s49_i),
.s50_r(s50_r),
.s50_i(s50_i),
.s51_r(s51_r),
.s51_i(s51_i),
.s52_r(s52_r),
.s52_i(s52_i),
.s53_r(s53_r),
.s53_i(s53_i),
.s54_r(s54_r),
.s54_i(s54_i),
.s55_r(s55_r),
.s55_i(s55_i),
.s56_r(s56_r),
.s56_i(s56_i),
.s57_r(s57_r),
.s57_i(s57_i),
.s58_r(s58_r),
.s58_i(s58_i),
.s59_r(s59_r),
.s59_i(s59_i),
.s60_r(s60_r),
.s60_i(s60_i),
.s61_r(s61_r),
.s61_i(s61_i),
.s62_r(s62_r),
.s62_i(s62_i),
.s63_r(s63_r),
.s63_i(s63_i),
.s64_r(s64_r),
.s64_i(s64_i),
.s65_r(s65_r),
.s65_i(s65_i),
.s66_r(s66_r),
.s66_i(s66_i),
.s67_r(s67_r),
.s67_i(s67_i),
.s68_r(s68_r),
.s68_i(s68_i),
.s69_r(s69_r),
.s69_i(s69_i),
.s70_r(s70_r),
.s70_i(s70_i),
.s71_r(s71_r),
.s71_i(s71_i),
.s72_r(s72_r),
.s72_i(s72_i),
.s73_r(s73_r),
.s73_i(s73_i),
.s74_r(s74_r),
.s74_i(s74_i),
.s75_r(s75_r),
.s75_i(s75_i),
.s76_r(s76_r),
.s76_i(s76_i),
.s77_r(s77_r),
.s77_i(s77_i),
.s78_r(s78_r),
.s78_i(s78_i),
.s79_r(s79_r),
.s79_i(s79_i),
.s80_r(s80_r),
.s80_i(s80_i),
.s81_r(s81_r),
.s81_i(s81_i),
.s82_r(s82_r),
.s82_i(s82_i),
.s83_r(s83_r),
.s83_i(s83_i),
.s84_r(s84_r),
.s84_i(s84_i),
.s85_r(s85_r),
.s85_i(s85_i),
.s86_r(s86_r),
.s86_i(s86_i),
.s87_r(s87_r),
.s87_i(s87_i),
.s88_r(s88_r),
.s88_i(s88_i),
.s89_r(s89_r),
.s89_i(s89_i),
.s90_r(s90_r),
.s90_i(s90_i),
.s91_r(s91_r),
.s91_i(s91_i),
.s92_r(s92_r),
.s92_i(s92_i),
.s93_r(s93_r),
.s93_i(s93_i),
.s94_r(s94_r),
.s94_i(s94_i),
.s95_r(s95_r),
.s95_i(s95_i),
.s96_r(s96_r),
.s96_i(s96_i),
.s97_r(s97_r),
.s97_i(s97_i),
.s98_r(s98_r),
.s98_i(s98_i),
.s99_r(s99_r),
.s99_i(s99_i),
.s100_r(s100_r),
.s100_i(s100_i),
.s101_r(s101_r),
.s101_i(s101_i),
.s102_r(s102_r),
.s102_i(s102_i),
.s103_r(s103_r),
.s103_i(s103_i),
.s104_r(s104_r),
.s104_i(s104_i),
.s105_r(s105_r),
.s105_i(s105_i),
.s106_r(s106_r),
.s106_i(s106_i),
.s107_r(s107_r),
.s107_i(s107_i),
.s108_r(s108_r),
.s108_i(s108_i),
.s109_r(s109_r),
.s109_i(s109_i),
.s110_r(s110_r),
.s110_i(s110_i),
.s111_r(s111_r),
.s111_i(s111_i),
.s112_r(s112_r),
.s112_i(s112_i),
.s113_r(s113_r),
.s113_i(s113_i),
.s114_r(s114_r),
.s114_i(s114_i),
.s115_r(s115_r),
.s115_i(s115_i),
.s116_r(s116_r),
.s116_i(s116_i),
.s117_r(s117_r),
.s117_i(s117_i),
.s118_r(s118_r),
.s118_i(s118_i),
.s119_r(s119_r),
.s119_i(s119_i),
.s120_r(s120_r),
.s120_i(s120_i),
.s121_r(s121_r),
.s121_i(s121_i),
.s122_r(s122_r),
.s122_i(s122_i),
.s123_r(s123_r),
.s123_i(s123_i),
.s124_r(s124_r),
.s124_i(s124_i),
.s125_r(s125_r),
.s125_i(s125_i),
.s126_r(s126_r),
.s126_i(s126_i),
.s127_r(s127_r),
.s127_i(s127_i),






.twiddle1_r(out_reg_twiddle_r_0),
.twiddle2_r(out_reg_twiddle_r_1),
.twiddle3_r(out_reg_twiddle_r_2),
.twiddle4_r(out_reg_twiddle_r_3),
.twiddle5_r(out_reg_twiddle_r_4),
.twiddle6_r(out_reg_twiddle_r_5),
.twiddle7_r(out_reg_twiddle_r_6),
.twiddle8_r(out_reg_twiddle_r_7),
.twiddle9_r(out_reg_twiddle_r_8),
.twiddle10_r(out_reg_twiddle_r_9),
.twiddle11_r(out_reg_twiddle_r_10),
.twiddle12_r(out_reg_twiddle_r_11),
.twiddle13_r(out_reg_twiddle_r_12),
.twiddle14_r(out_reg_twiddle_r_13),
.twiddle15_r(out_reg_twiddle_r_14),
.twiddle16_r(out_reg_twiddle_r_15),
.twiddle17_r(out_reg_twiddle_r_16),
.twiddle18_r(out_reg_twiddle_r_17),
.twiddle19_r(out_reg_twiddle_r_18),
.twiddle20_r(out_reg_twiddle_r_19),
.twiddle21_r(out_reg_twiddle_r_20),
.twiddle22_r(out_reg_twiddle_r_21),
.twiddle23_r(out_reg_twiddle_r_22),
.twiddle24_r(out_reg_twiddle_r_23),
.twiddle25_r(out_reg_twiddle_r_24),
.twiddle26_r(out_reg_twiddle_r_25),
.twiddle27_r(out_reg_twiddle_r_26),
.twiddle28_r(out_reg_twiddle_r_27),
.twiddle29_r(out_reg_twiddle_r_28),
.twiddle30_r(out_reg_twiddle_r_29),
.twiddle31_r(out_reg_twiddle_r_30),
.twiddle32_r(out_reg_twiddle_r_31),
.twiddle33_r(out_reg_twiddle_r_32),
.twiddle34_r(out_reg_twiddle_r_33),
.twiddle35_r(out_reg_twiddle_r_34),
.twiddle36_r(out_reg_twiddle_r_35),
.twiddle37_r(out_reg_twiddle_r_36),
.twiddle38_r(out_reg_twiddle_r_37),
.twiddle39_r(out_reg_twiddle_r_38),
.twiddle40_r(out_reg_twiddle_r_39),
.twiddle41_r(out_reg_twiddle_r_40),
.twiddle42_r(out_reg_twiddle_r_41),
.twiddle43_r(out_reg_twiddle_r_42),
.twiddle44_r(out_reg_twiddle_r_43),
.twiddle45_r(out_reg_twiddle_r_44),
.twiddle46_r(out_reg_twiddle_r_45),
.twiddle47_r(out_reg_twiddle_r_46),
.twiddle48_r(out_reg_twiddle_r_47),
.twiddle49_r(out_reg_twiddle_r_48),
.twiddle50_r(out_reg_twiddle_r_49),
.twiddle51_r(out_reg_twiddle_r_50),
.twiddle52_r(out_reg_twiddle_r_51),
.twiddle53_r(out_reg_twiddle_r_52),
.twiddle54_r(out_reg_twiddle_r_53),
.twiddle55_r(out_reg_twiddle_r_54),
.twiddle56_r(out_reg_twiddle_r_55),
.twiddle57_r(out_reg_twiddle_r_56),
.twiddle58_r(out_reg_twiddle_r_57),
.twiddle59_r(out_reg_twiddle_r_58),
.twiddle60_r(out_reg_twiddle_r_59),
.twiddle61_r(out_reg_twiddle_r_60),
.twiddle62_r(out_reg_twiddle_r_61),
.twiddle63_r(out_reg_twiddle_r_62),
.twiddle64_r(out_reg_twiddle_r_63),



.twiddle1_i(out_reg_twiddle_i_0),
.twiddle2_i(out_reg_twiddle_i_1),
.twiddle3_i(out_reg_twiddle_i_2),
.twiddle4_i(out_reg_twiddle_i_3),
.twiddle5_i(out_reg_twiddle_i_4),
.twiddle6_i(out_reg_twiddle_i_5),
.twiddle7_i(out_reg_twiddle_i_6),
.twiddle8_i(out_reg_twiddle_i_7),
.twiddle9_i(out_reg_twiddle_i_8),
.twiddle10_i(out_reg_twiddle_i_9),
.twiddle11_i(out_reg_twiddle_i_10),
.twiddle12_i(out_reg_twiddle_i_11),
.twiddle13_i(out_reg_twiddle_i_12),
.twiddle14_i(out_reg_twiddle_i_13),
.twiddle15_i(out_reg_twiddle_i_14),
.twiddle16_i(out_reg_twiddle_i_15),
.twiddle17_i(out_reg_twiddle_i_16),
.twiddle18_i(out_reg_twiddle_i_17),
.twiddle19_i(out_reg_twiddle_i_18),
.twiddle20_i(out_reg_twiddle_i_19),
.twiddle21_i(out_reg_twiddle_i_20),
.twiddle22_i(out_reg_twiddle_i_21),
.twiddle23_i(out_reg_twiddle_i_22),
.twiddle24_i(out_reg_twiddle_i_23),
.twiddle25_i(out_reg_twiddle_i_24),
.twiddle26_i(out_reg_twiddle_i_25),
.twiddle27_i(out_reg_twiddle_i_26),
.twiddle28_i(out_reg_twiddle_i_27),
.twiddle29_i(out_reg_twiddle_i_28),
.twiddle30_i(out_reg_twiddle_i_29),
.twiddle31_i(out_reg_twiddle_i_30),
.twiddle32_i(out_reg_twiddle_i_31),
.twiddle33_i(out_reg_twiddle_i_32),
.twiddle34_i(out_reg_twiddle_i_33),
.twiddle35_i(out_reg_twiddle_i_34),
.twiddle36_i(out_reg_twiddle_i_35),
.twiddle37_i(out_reg_twiddle_i_36),
.twiddle38_i(out_reg_twiddle_i_37),
.twiddle39_i(out_reg_twiddle_i_38),
.twiddle40_i(out_reg_twiddle_i_39),
.twiddle41_i(out_reg_twiddle_i_40),
.twiddle42_i(out_reg_twiddle_i_41),
.twiddle43_i(out_reg_twiddle_i_42),
.twiddle44_i(out_reg_twiddle_i_43),
.twiddle45_i(out_reg_twiddle_i_44),
.twiddle46_i(out_reg_twiddle_i_45),
.twiddle47_i(out_reg_twiddle_i_46),
.twiddle48_i(out_reg_twiddle_i_47),
.twiddle49_i(out_reg_twiddle_i_48),
.twiddle50_i(out_reg_twiddle_i_49),
.twiddle51_i(out_reg_twiddle_i_50),
.twiddle52_i(out_reg_twiddle_i_51),
.twiddle53_i(out_reg_twiddle_i_52),
.twiddle54_i(out_reg_twiddle_i_53),
.twiddle55_i(out_reg_twiddle_i_54),
.twiddle56_i(out_reg_twiddle_i_55),
.twiddle57_i(out_reg_twiddle_i_56),
.twiddle58_i(out_reg_twiddle_i_57),
.twiddle59_i(out_reg_twiddle_i_58),
.twiddle60_i(out_reg_twiddle_i_59),
.twiddle61_i(out_reg_twiddle_i_60),
.twiddle62_i(out_reg_twiddle_i_61),
.twiddle63_i(out_reg_twiddle_i_62),
.twiddle64_i(out_reg_twiddle_i_63)


);



twiddle_ROM_real_0 unt0
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_0)
 );

twiddle_ROM_real_1 unt1
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_1)
 );

twiddle_ROM_real_2 unt2
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_2)
 );

twiddle_ROM_real_3 unt3
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_3)
 );

twiddle_ROM_real_4 unt4
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_4)
 );

twiddle_ROM_real_5 unt5
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_5)
 );

twiddle_ROM_real_6 unt6
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_6)
 );

twiddle_ROM_real_7 unt7
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_7)
 );

twiddle_ROM_real_8 unt8
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_8)
 );

twiddle_ROM_real_9 unt9
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_9)
 );

twiddle_ROM_real_10 unt10
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_10)
 );

twiddle_ROM_real_11 unt11
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_11)
 );

twiddle_ROM_real_12 unt12
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_12)
 );

twiddle_ROM_real_13 unt13
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_13)
 );

twiddle_ROM_real_14 unt14
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_14)
 );

twiddle_ROM_real_15 unt15
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_r_15)
);





FFT_twiddle_ROM_img_0 unt_0
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_0)
 );

FFT_twiddle_ROM_img_1 unt_1
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_1)
 );

FFT_twiddle_ROM_img_2 unt_2
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_2)
 );

FFT_twiddle_ROM_img_3 unt_3
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_3)
 );

FFT_twiddle_ROM_img_4 unt_4
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_4)
 );

FFT_twiddle_ROM_img_5 unt_5
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_5)
 );

FFT_twiddle_ROM_img_6 unt_6
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_6)
 );

FFT_twiddle_ROM_img_7 unt_7
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_7)
 );

FFT_twiddle_ROM_img_8 unt_8
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_8)
 );

FFT_twiddle_ROM_img_9 unt_9
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_9)
 );

FFT_twiddle_ROM_img_10 unt_10
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_10)
 );

FFT_twiddle_ROM_img_11 unt_11
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_11)
 );

FFT_twiddle_ROM_img_12 unt_12
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_12)
 );

FFT_twiddle_ROM_img_13 unt_13
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_13)
 );

FFT_twiddle_ROM_img_14 unt_14
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_14)
 );

FFT_twiddle_ROM_img_15 unt_15
(
    .clk(clk),
    .addr(ROM_addr),
    .data_out(ROM_out_twiddle_i_15)
);





Controller_FSM #(.BITS(BITS),.NUMBER_OF_ENABLE_BITS(NUMBER_OF_ENABLE_BITS),.NUMBER_OF_MEM(NUMBER_OF_MEM),.MUX_SEL_BITS(SEL_BITS),.ADDRESS_BITS(ADDRESS_BITS)) U_Controller (
.ready_inputs(ready_inputs),
.clk(clk),
.rst(rst),
.reg_en(reg_en),
.twiddle_reg_en(twiddle_reg_en),
.ROM_addr(ROM_addr),
.correct(correct),
.sel_output_mux_0(sel_output_mux_0),
.sel_output_mux_1(sel_output_mux_1), 
.sel_output_mux_2(sel_output_mux_2), 
.sel_output_mux_3(sel_output_mux_3), 
.sel_output_mux_4(sel_output_mux_4), 
.sel_output_mux_5(sel_output_mux_5), 
.sel_output_mux_6(sel_output_mux_6), 
.sel_output_mux_7(sel_output_mux_7), 
.sel_output_mux_8(sel_output_mux_8), 
.sel_output_mux_9(sel_output_mux_9), 
.sel_output_mux_10(sel_output_mux_10), 
.sel_output_mux_11(sel_output_mux_11), 
.sel_output_mux_12(sel_output_mux_12), 
.sel_output_mux_13(sel_output_mux_13), 
.sel_output_mux_14(sel_output_mux_14), 
.sel_output_mux_15(sel_output_mux_15), 
.sel_output_mux_16(sel_output_mux_16), 
.sel_output_mux_17(sel_output_mux_17), 
.sel_output_mux_18(sel_output_mux_18), 
.sel_output_mux_19(sel_output_mux_19), 
.sel_output_mux_20(sel_output_mux_20), 
.sel_output_mux_21(sel_output_mux_21), 
.sel_output_mux_22(sel_output_mux_22), 
.sel_output_mux_23(sel_output_mux_23), 
.sel_output_mux_24(sel_output_mux_24), 
.sel_output_mux_25(sel_output_mux_25), 
.sel_output_mux_26(sel_output_mux_26), 
.sel_output_mux_27(sel_output_mux_27), 
.sel_output_mux_28(sel_output_mux_28), 
.sel_output_mux_29(sel_output_mux_29), 
.sel_output_mux_30(sel_output_mux_30), 
.sel_output_mux_31(sel_output_mux_31),
.read_address(read_address),
.write_address(write_address),
.mem_write_enable(mem_write_enable),
.sel_mux_2_1(sel_mux_2_1),
.sel_output_4x1 (sel_output_4x1)
);

MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U0_MUX_REAL_MEMORY (
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_0),
.mux_output(mux_0_output_real)
);

MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U1_MUX_REAL_MEMORY (
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_1),
.mux_output(mux_1_output_real)
);

MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U2_MUX_REAL_MEMORY (
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_2),
.mux_output(mux_2_output_real)
);

 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U3_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_3),
.mux_output(mux_3_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U4_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_4),
.mux_output(mux_4_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U5_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_5),
.mux_output(mux_5_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U6_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_6),
.mux_output(mux_6_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U7_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_7),
.mux_output(mux_7_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U8_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_8),
.mux_output(mux_8_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U9_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_9),
.mux_output(mux_9_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U10_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_10),
.mux_output(mux_10_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U11_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_11),
.mux_output(mux_11_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U12_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_12),
.mux_output(mux_12_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U13_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_13),
.mux_output(mux_13_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U14_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_14),
.mux_output(mux_14_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U15_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 

.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_15),
.mux_output(mux_15_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U16_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_16),
.mux_output(mux_16_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U17_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_17),
.mux_output(mux_17_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U18_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_18),
.mux_output(mux_18_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U19_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_19),
.mux_output(mux_19_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U20_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_20),
.mux_output(mux_20_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U21_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 

.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_21),
.mux_output(mux_21_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U22_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_22),
.mux_output(mux_22_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U23_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_23),
.mux_output(mux_23_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U24_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_24),
.mux_output(mux_24_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U25_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_25),
.mux_output(mux_25_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U26_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_26),
.mux_output(mux_26_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U27_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_27),
.mux_output(mux_27_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U28_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_28),
.mux_output(mux_28_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U29_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_29),
.mux_output(mux_29_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U30_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_30),
.mux_output(mux_30_output_real)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U31_MUX_REAL_MEMORY ( 
.mux_input_0(s0_r) , 
.mux_input_1(s1_r) , 
.mux_input_2(s2_r) , 
.mux_input_3(s3_r) , 
.mux_input_4(s4_r) , 
.mux_input_5(s5_r) , 
.mux_input_6(s6_r) , 
.mux_input_7(s7_r) , 
.mux_input_8(s8_r) , 
.mux_input_9(s9_r) , 
.mux_input_10(s10_r) , 
.mux_input_11(s11_r) , 
.mux_input_12(s12_r) , 
.mux_input_13(s13_r) , 
.mux_input_14(s14_r) , 
.mux_input_15(s15_r) , 
.mux_input_16(s16_r) , 
.mux_input_17(s17_r) , 
.mux_input_18(s18_r) , 
.mux_input_19(s19_r) , 
.mux_input_20(s20_r) , 
.mux_input_21(s21_r) , 
.mux_input_22(s22_r) , 
.mux_input_23(s23_r) , 
.mux_input_24(s24_r) , 
.mux_input_25(s25_r) , 
.mux_input_26(s26_r) , 
.mux_input_27(s27_r) , 
.mux_input_28(s28_r) , 
.mux_input_29(s29_r) , 
.mux_input_30(s30_r) , 
.mux_input_31(s31_r) , 
.mux_input_32(s32_r) , 
.mux_input_33(s33_r) , 
.mux_input_34(s34_r) , 
.mux_input_35(s35_r) , 
.mux_input_36(s36_r) , 
.mux_input_37(s37_r) , 
.mux_input_38(s38_r) , 
.mux_input_39(s39_r) , 
.mux_input_40(s40_r) , 
.mux_input_41(s41_r) , 
.mux_input_42(s42_r) , 
.mux_input_43(s43_r) , 
.mux_input_44(s44_r) , 
.mux_input_45(s45_r) , 
.mux_input_46(s46_r) , 
.mux_input_47(s47_r) , 
.mux_input_48(s48_r) , 
.mux_input_49(s49_r) , 
.mux_input_50(s50_r) , 
.mux_input_51(s51_r) , 
.mux_input_52(s52_r) , 
.mux_input_53(s53_r) , 
.mux_input_54(s54_r) , 
.mux_input_55(s55_r) , 
.mux_input_56(s56_r) , 
.mux_input_57(s57_r) , 
.mux_input_58(s58_r) , 
.mux_input_59(s59_r) , 
.mux_input_60(s60_r) , 
.mux_input_61(s61_r) , 
.mux_input_62(s62_r) , 
.mux_input_63(s63_r) , 
.mux_input_64(s64_r) , 
.mux_input_65(s65_r) , 
.mux_input_66(s66_r) , 
.mux_input_67(s67_r) , 
.mux_input_68(s68_r) , 
.mux_input_69(s69_r) , 
.mux_input_70(s70_r) , 
.mux_input_71(s71_r) , 
.mux_input_72(s72_r) , 
.mux_input_73(s73_r) , 
.mux_input_74(s74_r) , 
.mux_input_75(s75_r) , 
.mux_input_76(s76_r) , 
.mux_input_77(s77_r) , 
.mux_input_78(s78_r) , 
.mux_input_79(s79_r) , 
.mux_input_80(s80_r) , 
.mux_input_81(s81_r) , 
.mux_input_82(s82_r) , 
.mux_input_83(s83_r) , 
.mux_input_84(s84_r) , 
.mux_input_85(s85_r) , 
.mux_input_86(s86_r) , 
.mux_input_87(s87_r) , 
.mux_input_88(s88_r) , 
.mux_input_89(s89_r) , 
.mux_input_90(s90_r) , 
.mux_input_91(s91_r) , 
.mux_input_92(s92_r) , 
.mux_input_93(s93_r) , 
.mux_input_94(s94_r) , 
.mux_input_95(s95_r) , 
.mux_input_96(s96_r) , 
.mux_input_97(s97_r) , 
.mux_input_98(s98_r) , 
.mux_input_99(s99_r) , 
.mux_input_100(s100_r) , 
.mux_input_101(s101_r) , 
.mux_input_102(s102_r) , 
.mux_input_103(s103_r) , 
.mux_input_104(s104_r) , 
.mux_input_105(s105_r) , 
.mux_input_106(s106_r) , 
.mux_input_107(s107_r) , 
.mux_input_108(s108_r) , 
.mux_input_109(s109_r) , 
.mux_input_110(s110_r) , 
.mux_input_111(s111_r) , 
.mux_input_112(s112_r) , 
.mux_input_113(s113_r) , 
.mux_input_114(s114_r) , 
.mux_input_115(s115_r) , 
.mux_input_116(s116_r) , 
.mux_input_117(s117_r) , 
.mux_input_118(s118_r) , 
.mux_input_119(s119_r) , 
.mux_input_120(s120_r) , 
.mux_input_121(s121_r) , 
.mux_input_122(s122_r) , 
.mux_input_123(s123_r) , 
.mux_input_124(s124_r) , 
.mux_input_125(s125_r) , 
.mux_input_126(s126_r) , 
.mux_input_127(s127_r) ,
.sel_input(sel_output_mux_31),
.mux_output(mux_31_output_real));

MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U0_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_0),
.mux_output(mux_0_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U1_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_1),
.mux_output(mux_1_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U2_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_2),
.mux_output(mux_2_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U3_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_3),
.mux_output(mux_3_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U4_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_4),
.mux_output(mux_4_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U5_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_5),
.mux_output(mux_5_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U6_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_6),
.mux_output(mux_6_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U7_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_7),
.mux_output(mux_7_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U8_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_8),
.mux_output(mux_8_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U9_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_9),
.mux_output(mux_9_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U10_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_10),
.mux_output(mux_10_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U11_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_11),
.mux_output(mux_11_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U12_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_12),
.mux_output(mux_12_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U13_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_13),
.mux_output(mux_13_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U14_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_14),
.mux_output(mux_14_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U15_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_15),
.mux_output(mux_15_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U16_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_16),
.mux_output(mux_16_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U17_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_17),
.mux_output(mux_17_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U18_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_18),
.mux_output(mux_18_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U19_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_19),
.mux_output(mux_19_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U20_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_20),
.mux_output(mux_20_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U21_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_21),
.mux_output(mux_21_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U22_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_22),
.mux_output(mux_22_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U23_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_23),
.mux_output(mux_23_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U24_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_24),
.mux_output(mux_24_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U25_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_25),
.mux_output(mux_25_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U26_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_26),
.mux_output(mux_26_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U27_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_27),
.mux_output(mux_27_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U28_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_28),
.mux_output(mux_28_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U29_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_29),
.mux_output(mux_29_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U30_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_30),
.mux_output(mux_30_output_imag)); 
 
MUX_128_1 #(.BITS(BITS),.SEL_BITS(SEL_BITS)) U31_MUX_IMAG_MEMORY ( 
.mux_input_0(s0_i) , 
.mux_input_1(s1_i) , 
.mux_input_2(s2_i) , 
.mux_input_3(s3_i) , 
.mux_input_4(s4_i) , 
.mux_input_5(s5_i) , 
.mux_input_6(s6_i) , 
.mux_input_7(s7_i) , 
.mux_input_8(s8_i) , 
.mux_input_9(s9_i) , 
.mux_input_10(s10_i) , 
.mux_input_11(s11_i) , 
.mux_input_12(s12_i) , 
.mux_input_13(s13_i) , 
.mux_input_14(s14_i) , 
.mux_input_15(s15_i) , 
.mux_input_16(s16_i) , 
.mux_input_17(s17_i) , 
.mux_input_18(s18_i) , 
.mux_input_19(s19_i) , 
.mux_input_20(s20_i) , 
.mux_input_21(s21_i) , 
.mux_input_22(s22_i) , 
.mux_input_23(s23_i) , 
.mux_input_24(s24_i) , 
.mux_input_25(s25_i) , 
.mux_input_26(s26_i) , 
.mux_input_27(s27_i) , 
.mux_input_28(s28_i) , 
.mux_input_29(s29_i) , 
.mux_input_30(s30_i) , 
.mux_input_31(s31_i) , 
.mux_input_32(s32_i) , 
.mux_input_33(s33_i) , 
.mux_input_34(s34_i) , 
.mux_input_35(s35_i) , 
.mux_input_36(s36_i) , 
.mux_input_37(s37_i) , 
.mux_input_38(s38_i) , 
.mux_input_39(s39_i) , 
.mux_input_40(s40_i) , 
.mux_input_41(s41_i) , 
.mux_input_42(s42_i) , 
.mux_input_43(s43_i) , 
.mux_input_44(s44_i) , 
.mux_input_45(s45_i) , 
.mux_input_46(s46_i) , 
.mux_input_47(s47_i) , 
.mux_input_48(s48_i) , 
.mux_input_49(s49_i) , 
.mux_input_50(s50_i) , 
.mux_input_51(s51_i) , 
.mux_input_52(s52_i) , 
.mux_input_53(s53_i) , 
.mux_input_54(s54_i) , 
.mux_input_55(s55_i) , 
.mux_input_56(s56_i) , 
.mux_input_57(s57_i) , 
.mux_input_58(s58_i) , 
.mux_input_59(s59_i) , 
.mux_input_60(s60_i) , 
.mux_input_61(s61_i) , 
.mux_input_62(s62_i) , 
.mux_input_63(s63_i) , 
.mux_input_64(s64_i) , 
.mux_input_65(s65_i) , 
.mux_input_66(s66_i) , 
.mux_input_67(s67_i) , 
.mux_input_68(s68_i) , 
.mux_input_69(s69_i) , 
.mux_input_70(s70_i) , 
.mux_input_71(s71_i) , 
.mux_input_72(s72_i) , 
.mux_input_73(s73_i) , 
.mux_input_74(s74_i) , 
.mux_input_75(s75_i) , 
.mux_input_76(s76_i) , 
.mux_input_77(s77_i) , 
.mux_input_78(s78_i) , 
.mux_input_79(s79_i) , 
.mux_input_80(s80_i) , 
.mux_input_81(s81_i) , 
.mux_input_82(s82_i) , 
.mux_input_83(s83_i) , 
.mux_input_84(s84_i) , 
.mux_input_85(s85_i) , 
.mux_input_86(s86_i) , 
.mux_input_87(s87_i) , 
.mux_input_88(s88_i) , 
.mux_input_89(s89_i) , 
.mux_input_90(s90_i) , 
.mux_input_91(s91_i) , 
.mux_input_92(s92_i) , 
.mux_input_93(s93_i) , 
.mux_input_94(s94_i) , 
.mux_input_95(s95_i) , 
.mux_input_96(s96_i) , 
.mux_input_97(s97_i) , 
.mux_input_98(s98_i) , 
.mux_input_99(s99_i) , 
.mux_input_100(s100_i) , 
.mux_input_101(s101_i) , 
.mux_input_102(s102_i) , 
.mux_input_103(s103_i) , 
.mux_input_104(s104_i) , 
.mux_input_105(s105_i) , 
.mux_input_106(s106_i) , 
.mux_input_107(s107_i) , 
.mux_input_108(s108_i) , 
.mux_input_109(s109_i) , 
.mux_input_110(s110_i) , 
.mux_input_111(s111_i) , 
.mux_input_112(s112_i) , 
.mux_input_113(s113_i) , 
.mux_input_114(s114_i) , 
.mux_input_115(s115_i) , 
.mux_input_116(s116_i) , 
.mux_input_117(s117_i) , 
.mux_input_118(s118_i) , 
.mux_input_119(s119_i) , 
.mux_input_120(s120_i) , 
.mux_input_121(s121_i) , 
.mux_input_122(s122_i) , 
.mux_input_123(s123_i) , 
.mux_input_124(s124_i) , 
.mux_input_125(s125_i) , 
.mux_input_126(s126_i) , 
.mux_input_127(s127_i) ,
.sel_input(sel_output_mux_31),
.mux_output(mux_31_output_imag)); 
 

Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U0_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_0_output_real),
.write_enable(mem_write_enable[0]),
.read_data(memory_real_output_0));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U1_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_1_output_real),
.write_enable(mem_write_enable[1]),
.read_data(memory_real_output_1));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U2_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_2_output_real),
.write_enable(mem_write_enable[2]),
.read_data(memory_real_output_2));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U3_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_3_output_real),
.write_enable(mem_write_enable[3]),
.read_data(memory_real_output_3));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U4_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_4_output_real),
.write_enable(mem_write_enable[4]),
.read_data(memory_real_output_4));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U5_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_5_output_real),
.write_enable(mem_write_enable[5]),
.read_data(memory_real_output_5));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U6_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_6_output_real),
.write_enable(mem_write_enable[6]),
.read_data(memory_real_output_6));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U7_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_7_output_real),
.write_enable(mem_write_enable[7]),
.read_data(memory_real_output_7));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U8_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_8_output_real),
.write_enable(mem_write_enable[8]),
.read_data(memory_real_output_8));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U9_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_9_output_real),
.write_enable(mem_write_enable[9]),
.read_data(memory_real_output_9));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U10_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_10_output_real),
.write_enable(mem_write_enable[10]),
.read_data(memory_real_output_10));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U11_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_11_output_real),
.write_enable(mem_write_enable[11]),
.read_data(memory_real_output_11));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U12_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_12_output_real),
.write_enable(mem_write_enable[12]),
.read_data(memory_real_output_12));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U13_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_13_output_real),
.write_enable(mem_write_enable[13]),
.read_data(memory_real_output_13));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U14_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_14_output_real),
.write_enable(mem_write_enable[14]),
.read_data(memory_real_output_14));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U15_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_15_output_real),
.write_enable(mem_write_enable[15]),
.read_data(memory_real_output_15));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U16_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_16_output_real),
.write_enable(mem_write_enable[16]),
.read_data(memory_real_output_16));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U17_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_17_output_real),
.write_enable(mem_write_enable[17]),
.read_data(memory_real_output_17));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U18_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_18_output_real),
.write_enable(mem_write_enable[18]),
.read_data(memory_real_output_18));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U19_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_19_output_real),
.write_enable(mem_write_enable[19]),
.read_data(memory_real_output_19));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U20_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_20_output_real),
.write_enable(mem_write_enable[20]),
.read_data(memory_real_output_20));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U21_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_21_output_real),
.write_enable(mem_write_enable[21]),
.read_data(memory_real_output_21));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U22_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_22_output_real),
.write_enable(mem_write_enable[22]),
.read_data(memory_real_output_22));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U23_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_23_output_real),
.write_enable(mem_write_enable[23]),
.read_data(memory_real_output_23));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U24_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_24_output_real),
.write_enable(mem_write_enable[24]),
.read_data(memory_real_output_24));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U25_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_25_output_real),
.write_enable(mem_write_enable[25]),
.read_data(memory_real_output_25));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U26_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_26_output_real),
.write_enable(mem_write_enable[26]),
.read_data(memory_real_output_26));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U27_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_27_output_real),
.write_enable(mem_write_enable[27]),
.read_data(memory_real_output_27));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U28_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_28_output_real),
.write_enable(mem_write_enable[28]),
.read_data(memory_real_output_28));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U29_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_29_output_real),
.write_enable(mem_write_enable[29]),
.read_data(memory_real_output_29));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U30_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_30_output_real),
.write_enable(mem_write_enable[30]),
.read_data(memory_real_output_30));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U31_REAL_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_31_output_real),
.write_enable(mem_write_enable[31]),
.read_data(memory_real_output_31));
 

Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U0_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_0_output_imag),
.write_enable(mem_write_enable[0]),
.read_data(memory_imag_output_0));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U1_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_1_output_imag),
.write_enable(mem_write_enable[1]),
.read_data(memory_imag_output_1));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U2_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_2_output_imag),
.write_enable(mem_write_enable[2]),
.read_data(memory_imag_output_2));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U3_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_3_output_imag),
.write_enable(mem_write_enable[3]),
.read_data(memory_imag_output_3));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U4_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_4_output_imag),
.write_enable(mem_write_enable[4]),
.read_data(memory_imag_output_4));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U5_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_5_output_imag),
.write_enable(mem_write_enable[5]),
.read_data(memory_imag_output_5));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U6_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_6_output_imag),
.write_enable(mem_write_enable[6]),
.read_data(memory_imag_output_6));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U7_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_7_output_imag),
.write_enable(mem_write_enable[7]),
.read_data(memory_imag_output_7));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U8_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_8_output_imag),
.write_enable(mem_write_enable[8]),
.read_data(memory_imag_output_8));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U9_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_9_output_imag),
.write_enable(mem_write_enable[9]),
.read_data(memory_imag_output_9));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U10_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_10_output_imag),
.write_enable(mem_write_enable[10]),
.read_data(memory_imag_output_10));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U11_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_11_output_imag),
.write_enable(mem_write_enable[11]),
.read_data(memory_imag_output_11));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U12_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_12_output_imag),
.write_enable(mem_write_enable[12]),
.read_data(memory_imag_output_12));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U13_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_13_output_imag),
.write_enable(mem_write_enable[13]),
.read_data(memory_imag_output_13));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U14_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_14_output_imag),
.write_enable(mem_write_enable[14]),
.read_data(memory_imag_output_14));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U15_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_15_output_imag),
.write_enable(mem_write_enable[15]),
.read_data(memory_imag_output_15));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U16_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_16_output_imag),
.write_enable(mem_write_enable[16]),
.read_data(memory_imag_output_16));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U17_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_17_output_imag),
.write_enable(mem_write_enable[17]),
.read_data(memory_imag_output_17));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U18_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_18_output_imag),
.write_enable(mem_write_enable[18]),
.read_data(memory_imag_output_18));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U19_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_19_output_imag),
.write_enable(mem_write_enable[19]),
.read_data(memory_imag_output_19));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U20_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_20_output_imag),
.write_enable(mem_write_enable[20]),
.read_data(memory_imag_output_20));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U21_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_21_output_imag),
.write_enable(mem_write_enable[21]),
.read_data(memory_imag_output_21));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U22_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_22_output_imag),
.write_enable(mem_write_enable[22]),
.read_data(memory_imag_output_22));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U23_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_23_output_imag),
.write_enable(mem_write_enable[23]),
.read_data(memory_imag_output_23));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U24_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_24_output_imag),
.write_enable(mem_write_enable[24]),
.read_data(memory_imag_output_24));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U25_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_25_output_imag),
.write_enable(mem_write_enable[25]),
.read_data(memory_imag_output_25));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U26_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_26_output_imag),
.write_enable(mem_write_enable[26]),
.read_data(memory_imag_output_26));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U27_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_27_output_imag),
.write_enable(mem_write_enable[27]),
.read_data(memory_imag_output_27));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U28_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_28_output_imag),
.write_enable(mem_write_enable[28]),
.read_data(memory_imag_output_28));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U29_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_29_output_imag),
.write_enable(mem_write_enable[29]),
.read_data(memory_imag_output_29));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U30_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_30_output_imag),
.write_enable(mem_write_enable[30]),
.read_data(memory_imag_output_30));
 
Memory #(.BITS(BITS),.ADDRESS_BITS(ADDRESS_BITS),.NUMBER_OF_LOCATIONS(NUMBER_OF_LOCATIONS)) U31_IMAG_MEMORY (
.clk(clk),
.rst(rst),
.read_address(read_address),
.write_address(write_address),
.write_data(mux_2_1_31_output_imag),
.write_enable(mem_write_enable[31]),
.read_data(memory_imag_output_31));
 
MUX_2_1 #(.BITS(BITS)) U0_REAL_MUX_2_1 (
    .in_1(mux4_mux2_0_r),
    .in_2(mux_0_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_0_output_real)
);

MUX_2_1 #(.BITS(BITS)) U1_REAL_MUX_2_1 (
    .in_1(mux4_mux2_1_r),
    .in_2(mux_1_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_1_output_real)
);

MUX_2_1 #(.BITS(BITS)) U2_REAL_MUX_2_1 (
    .in_1(mux4_mux2_2_r),
    .in_2(mux_2_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_2_output_real)
);

MUX_2_1 #(.BITS(BITS)) U3_REAL_MUX_2_1 (
    .in_1(mux4_mux2_3_r),
    .in_2(mux_3_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_3_output_real)
);

MUX_2_1 #(.BITS(BITS)) U4_REAL_MUX_2_1 (
    .in_1(mux4_mux2_4_r),
    .in_2(mux_4_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_4_output_real)
);

MUX_2_1 #(.BITS(BITS)) U5_REAL_MUX_2_1 (
    .in_1(mux4_mux2_5_r),
    .in_2(mux_5_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_5_output_real)
);

MUX_2_1 #(.BITS(BITS)) U6_REAL_MUX_2_1 (
    .in_1(mux4_mux2_6_r),
    .in_2(mux_6_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_6_output_real)
);

MUX_2_1 #(.BITS(BITS)) U7_REAL_MUX_2_1 (
    .in_1(mux4_mux2_7_r),
    .in_2(mux_7_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_7_output_real)
);

MUX_2_1 #(.BITS(BITS)) U8_REAL_MUX_2_1 (
    .in_1(mux4_mux2_8_r),
    .in_2(mux_8_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_8_output_real)
);

MUX_2_1 #(.BITS(BITS)) U9_REAL_MUX_2_1 (
    .in_1(mux4_mux2_9_r),
    .in_2(mux_9_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_9_output_real)
);

MUX_2_1 #(.BITS(BITS)) U10_REAL_MUX_2_1 (
    .in_1(mux4_mux2_10_r),
    .in_2(mux_10_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_10_output_real)
);

MUX_2_1 #(.BITS(BITS)) U11_REAL_MUX_2_1 (
    .in_1(mux4_mux2_11_r),
    .in_2(mux_11_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_11_output_real)
);

MUX_2_1 #(.BITS(BITS)) U12_REAL_MUX_2_1 (
    .in_1(mux4_mux2_12_r),
    .in_2(mux_12_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_12_output_real)
);

MUX_2_1 #(.BITS(BITS)) U13_REAL_MUX_2_1 (
    .in_1(mux4_mux2_13_r),
    .in_2(mux_13_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_13_output_real)
);

MUX_2_1 #(.BITS(BITS)) U14_REAL_MUX_2_1 (
    .in_1(mux4_mux2_14_r),
    .in_2(mux_14_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_14_output_real)
);

MUX_2_1 #(.BITS(BITS)) U15_REAL_MUX_2_1 (
    .in_1(mux4_mux2_15_r),
    .in_2(mux_15_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_15_output_real)
);

MUX_2_1 #(.BITS(BITS)) U16_REAL_MUX_2_1 (
    .in_1(mux4_mux2_16_r),
    .in_2(mux_16_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_16_output_real)
);

MUX_2_1 #(.BITS(BITS)) U17_REAL_MUX_2_1 (
    .in_1(mux4_mux2_17_r),
    .in_2(mux_17_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_17_output_real)
);

MUX_2_1 #(.BITS(BITS)) U18_REAL_MUX_2_1 (
    .in_1(mux4_mux2_18_r),
    .in_2(mux_18_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_18_output_real)
);

MUX_2_1 #(.BITS(BITS)) U19_REAL_MUX_2_1 (
    .in_1(mux4_mux2_19_r),
    .in_2(mux_19_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_19_output_real)
);

MUX_2_1 #(.BITS(BITS)) U20_REAL_MUX_2_1 (
    .in_1(mux4_mux2_20_r),
    .in_2(mux_20_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_20_output_real)
);

MUX_2_1 #(.BITS(BITS)) U21_REAL_MUX_2_1 (
    .in_1(mux4_mux2_21_r),
    .in_2(mux_21_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_21_output_real)
);

MUX_2_1 #(.BITS(BITS)) U22_REAL_MUX_2_1 (
    .in_1(mux4_mux2_22_r),
    .in_2(mux_22_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_22_output_real)
);

MUX_2_1 #(.BITS(BITS)) U23_REAL_MUX_2_1 (
    .in_1(mux4_mux2_23_r),
    .in_2(mux_23_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_23_output_real)
);

MUX_2_1 #(.BITS(BITS)) U24_REAL_MUX_2_1 (
    .in_1(mux4_mux2_24_r),
    .in_2(mux_24_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_24_output_real)
);

MUX_2_1 #(.BITS(BITS)) U25_REAL_MUX_2_1 (
    .in_1(mux4_mux2_25_r),
    .in_2(mux_25_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_25_output_real)
);

MUX_2_1 #(.BITS(BITS)) U26_REAL_MUX_2_1 (
    .in_1(mux4_mux2_26_r),
    .in_2(mux_26_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_26_output_real)
);

MUX_2_1 #(.BITS(BITS)) U27_REAL_MUX_2_1 (
    .in_1(mux4_mux2_27_r),
    .in_2(mux_27_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_27_output_real)
);

MUX_2_1 #(.BITS(BITS)) U28_REAL_MUX_2_1 (
    .in_1(mux4_mux2_28_r),
    .in_2(mux_28_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_28_output_real)
);

MUX_2_1 #(.BITS(BITS)) U29_REAL_MUX_2_1 (
    .in_1(mux4_mux2_29_r),
    .in_2(mux_29_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_29_output_real)
);

MUX_2_1 #(.BITS(BITS)) U30_REAL_MUX_2_1 (
    .in_1(mux4_mux2_30_r),
    .in_2(mux_30_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_30_output_real)
);

MUX_2_1 #(.BITS(BITS)) U31_REAL_MUX_2_1 (
    .in_1(mux4_mux2_31_r),
    .in_2(mux_31_output_real),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_31_output_real)
);


MUX_2_1 #(.BITS(BITS)) U0_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_0_i),
    .in_2(mux_0_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_0_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U1_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_1_i),
    .in_2(mux_1_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_1_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U2_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_2_i),
    .in_2(mux_2_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_2_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U3_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_3_i),
    .in_2(mux_3_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_3_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U4_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_4_i),
    .in_2(mux_4_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_4_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U5_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_5_i),
    .in_2(mux_5_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_5_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U6_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_6_i),
    .in_2(mux_6_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_6_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U7_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_7_i),
    .in_2(mux_7_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_7_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U8_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_8_i),
    .in_2(mux_8_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_8_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U9_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_9_i),
    .in_2(mux_9_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_9_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U10_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_10_i),
    .in_2(mux_10_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_10_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U11_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_11_i),
    .in_2(mux_11_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_11_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U12_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_12_i),
    .in_2(mux_12_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_12_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U13_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_13_i),
    .in_2(mux_13_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_13_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U14_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_14_i),
    .in_2(mux_14_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_14_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U15_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_15_i),
    .in_2(mux_15_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_15_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U16_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_16_i),
    .in_2(mux_16_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_16_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U17_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_17_i),
    .in_2(mux_17_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_17_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U18_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_18_i),
    .in_2(mux_18_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_18_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U19_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_19_i),
    .in_2(mux_19_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_19_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U20_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_20_i),
    .in_2(mux_20_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_20_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U21_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_21_i),
    .in_2(mux_21_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_21_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U22_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_22_i),
    .in_2(mux_22_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_22_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U23_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_23_i),
    .in_2(mux_23_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_23_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U24_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_24_i),
    .in_2(mux_24_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_24_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U25_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_25_i),
    .in_2(mux_25_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_25_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U26_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_26_i),
    .in_2(mux_26_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_26_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U27_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_27_i),
    .in_2(mux_27_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_27_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U28_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_28_i),
    .in_2(mux_28_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_28_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U29_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_29_i),
    .in_2(mux_29_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_29_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U30_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_30_i),
    .in_2(mux_30_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_30_output_imag)
);

MUX_2_1 #(.BITS(BITS)) U31_IMAG_MUX_2_1 (
    .in_1(mux4_mux2_31_i),
    .in_2(mux_31_output_imag),
    .selection_line(sel_mux_2_1),
    .out(mux_2_1_31_output_imag)
);




MUX_4_1 #(.BITS(BITS)) U0_MUX_REAL_4_1
(
    .in_0(x0_r),
    .in_1(x64_r),
    .in_2(x32_r),
    .in_3(x96_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_0_r)
);

MUX_4_1 #(.BITS(BITS)) U1_MUX_REAL_4_1
(
    .in_0(x16_r),
    .in_1(x80_r),
    .in_2(x48_r),
    .in_3(x112_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_1_r)
);

MUX_4_1 #(.BITS(BITS)) U2_MUX_REAL_4_1
(
    .in_0(x8_r),
    .in_1(x72_r),
    .in_2(x40_r),
    .in_3(x104_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_2_r)
);

MUX_4_1 #(.BITS(BITS)) U3_MUX_REAL_4_1
(
    .in_0(x24_r),
    .in_1(x88_r),
    .in_2(x56_r),
    .in_3(x120_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_3_r)
);

MUX_4_1 #(.BITS(BITS)) U4_MUX_REAL_4_1
(
    .in_0(x4_r),
    .in_1(x68_r),
    .in_2(x36_r),
    .in_3(x100_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_4_r)
);

MUX_4_1 #(.BITS(BITS)) U5_MUX_REAL_4_1
(
    .in_0(x20_r),
    .in_1(x84_r),
    .in_2(x52_r),
    .in_3(x116_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_5_r)
);

MUX_4_1 #(.BITS(BITS)) U6_MUX_REAL_4_1
(
    .in_0(x12_r),
    .in_1(x76_r),
    .in_2(x44_r),
    .in_3(x108_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_6_r)
);

MUX_4_1 #(.BITS(BITS)) U7_MUX_REAL_4_1
(
    .in_0(x28_r),
    .in_1(x92_r),
    .in_2(x60_r),
    .in_3(x124_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_7_r)
);

MUX_4_1 #(.BITS(BITS)) U8_MUX_REAL_4_1
(
    .in_0(x2_r),
    .in_1(x66_r),
    .in_2(x34_r),
    .in_3(x98_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_8_r)
);

MUX_4_1 #(.BITS(BITS)) U9_MUX_REAL_4_1
(
    .in_0(x18_r),
    .in_1(x82_r),
    .in_2(x50_r),
    .in_3(x114_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_9_r)
);

MUX_4_1 #(.BITS(BITS)) U10_MUX_REAL_4_1
(
    .in_0(x10_r),
    .in_1(x74_r),
    .in_2(x42_r),
    .in_3(x106_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_10_r)
);

MUX_4_1 #(.BITS(BITS)) U11_MUX_REAL_4_1
(
    .in_0(x26_r),
    .in_1(x90_r),
    .in_2(x58_r),
    .in_3(x122_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_11_r)
);

MUX_4_1 #(.BITS(BITS)) U12_MUX_REAL_4_1
(
    .in_0(x6_r),
    .in_1(x70_r),
    .in_2(x38_r),
    .in_3(x102_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_12_r)
);

MUX_4_1 #(.BITS(BITS)) U13_MUX_REAL_4_1
(
    .in_0(x22_r),
    .in_1(x86_r),
    .in_2(x54_r),
    .in_3(x118_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_13_r)
);

MUX_4_1 #(.BITS(BITS)) U14_MUX_REAL_4_1
(
    .in_0(x14_r),
    .in_1(x78_r),
    .in_2(x46_r),
    .in_3(x110_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_14_r)
);

MUX_4_1 #(.BITS(BITS)) U15_MUX_REAL_4_1
(
    .in_0(x30_r),
    .in_1(x94_r),
    .in_2(x62_r),
    .in_3(x126_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_15_r)
);

MUX_4_1 #(.BITS(BITS)) U16_MUX_REAL_4_1
(
    .in_0(x1_r),
    .in_1(x65_r),
    .in_2(x33_r),
    .in_3(x97_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_16_r)
);

MUX_4_1 #(.BITS(BITS)) U17_MUX_REAL_4_1
(
    .in_0(x17_r),
    .in_1(x81_r),
    .in_2(x49_r),
    .in_3(x113_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_17_r)
);

MUX_4_1 #(.BITS(BITS)) U18_MUX_REAL_4_1
(
    .in_0(x9_r),
    .in_1(x73_r),
    .in_2(x41_r),
    .in_3(x105_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_18_r)
);

MUX_4_1 #(.BITS(BITS)) U19_MUX_REAL_4_1
(
    .in_0(x25_r),
    .in_1(x89_r),
    .in_2(x57_r),
    .in_3(x121_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_19_r)
);

MUX_4_1 #(.BITS(BITS)) U20_MUX_REAL_4_1
(
    .in_0(x5_r),
    .in_1(x69_r),
    .in_2(x37_r),
    .in_3(x101_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_20_r)
);

MUX_4_1 #(.BITS(BITS)) U21_MUX_REAL_4_1
(
    .in_0(x21_r),
    .in_1(x85_r),
    .in_2(x53_r),
    .in_3(x117_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_21_r)
);

MUX_4_1 #(.BITS(BITS)) U22_MUX_REAL_4_1
(
    .in_0(x13_r),
    .in_1(x77_r),
    .in_2(x45_r),
    .in_3(x109_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_22_r)
);

MUX_4_1 #(.BITS(BITS)) U23_MUX_REAL_4_1
(
    .in_0(x29_r),
    .in_1(x93_r),
    .in_2(x61_r),
    .in_3(x125_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_23_r)
);

MUX_4_1 #(.BITS(BITS)) U24_MUX_REAL_4_1
(
    .in_0(x3_r),
    .in_1(x67_r),
    .in_2(x35_r),
    .in_3(x99_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_24_r)
);

MUX_4_1 #(.BITS(BITS)) U25_MUX_REAL_4_1
(
    .in_0(x19_r),
    .in_1(x83_r),
    .in_2(x51_r),
    .in_3(x115_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_25_r)
);

MUX_4_1 #(.BITS(BITS)) U26_MUX_REAL_4_1
(
    .in_0(x11_r),
    .in_1(x75_r),
    .in_2(x43_r),
    .in_3(x107_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_26_r)
);

MUX_4_1 #(.BITS(BITS)) U27_MUX_REAL_4_1
(
    .in_0(x27_r),
    .in_1(x91_r),
    .in_2(x59_r),
    .in_3(x123_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_27_r)
);

MUX_4_1 #(.BITS(BITS)) U28_MUX_REAL_4_1
(
    .in_0(x7_r),
    .in_1(x71_r),
    .in_2(x39_r),
    .in_3(x103_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_28_r)
);

MUX_4_1 #(.BITS(BITS)) U29_MUX_REAL_4_1
(
    .in_0(x23_r),
    .in_1(x87_r),
    .in_2(x55_r),
    .in_3(x119_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_29_r)
);

MUX_4_1 #(.BITS(BITS)) U30_MUX_REAL_4_1
(
    .in_0(x15_r),
    .in_1(x79_r),
    .in_2(x47_r),
    .in_3(x111_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_30_r)
);

MUX_4_1 #(.BITS(BITS)) U31_MUX_REAL_4_1
(
    .in_0(x31_r),
    .in_1(x95_r),
    .in_2(x63_r),
    .in_3(x127_r),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_31_r)
);



MUX_4_1 #(.BITS(BITS)) U0_MUX_IMAG_4_1
(
    .in_0(x0_i),
    .in_1(x64_i),
    .in_2(x32_i),
    .in_3(x96_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_0_i)
);

MUX_4_1 #(.BITS(BITS)) U1_MUX_IMAG_4_1
(
    .in_0(x16_i),
    .in_1(x80_i),
    .in_2(x48_i),
    .in_3(x112_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_1_i)
);

MUX_4_1 #(.BITS(BITS)) U2_MUX_IMAG_4_1
(
    .in_0(x8_i),
    .in_1(x72_i),
    .in_2(x40_i),
    .in_3(x104_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_2_i)
);

MUX_4_1 #(.BITS(BITS)) U3_MUX_IMAG_4_1
(
    .in_0(x24_i),
    .in_1(x88_i),
    .in_2(x56_i),
    .in_3(x120_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_3_i)
);

MUX_4_1 #(.BITS(BITS)) U4_MUX_IMAG_4_1
(
    .in_0(x4_i),
    .in_1(x68_i),
    .in_2(x36_i),
    .in_3(x100_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_4_i)
);

MUX_4_1 #(.BITS(BITS)) U5_MUX_IMAG_4_1
(
    .in_0(x20_i),
    .in_1(x84_i),
    .in_2(x52_i),
    .in_3(x116_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_5_i)
);

MUX_4_1 #(.BITS(BITS)) U6_MUX_IMAG_4_1
(
    .in_0(x12_i),
    .in_1(x76_i),
    .in_2(x44_i),
    .in_3(x108_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_6_i)
);

MUX_4_1 #(.BITS(BITS)) U7_MUX_IMAG_4_1
(
    .in_0(x28_i),
    .in_1(x92_i),
    .in_2(x60_i),
    .in_3(x124_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_7_i)
);

MUX_4_1 #(.BITS(BITS)) U8_MUX_IMAG_4_1
(
    .in_0(x2_i),
    .in_1(x66_i),
    .in_2(x34_i),
    .in_3(x98_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_8_i)
);

MUX_4_1 #(.BITS(BITS)) U9_MUX_IMAG_4_1
(
    .in_0(x18_i),
    .in_1(x82_i),
    .in_2(x50_i),
    .in_3(x114_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_9_i)
);

MUX_4_1 #(.BITS(BITS)) U10_MUX_IMAG_4_1
(
    .in_0(x10_i),
    .in_1(x74_i),
    .in_2(x42_i),
    .in_3(x106_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_10_i)
);

MUX_4_1 #(.BITS(BITS)) U11_MUX_IMAG_4_1
(
    .in_0(x26_i),
    .in_1(x90_i),
    .in_2(x58_i),
    .in_3(x122_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_11_i)
);

MUX_4_1 #(.BITS(BITS)) U12_MUX_IMAG_4_1
(
    .in_0(x6_i),
    .in_1(x70_i),
    .in_2(x38_i),
    .in_3(x102_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_12_i)
);

MUX_4_1 #(.BITS(BITS)) U13_MUX_IMAG_4_1
(
    .in_0(x22_i),
    .in_1(x86_i),
    .in_2(x54_i),
    .in_3(x118_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_13_i)
);

MUX_4_1 #(.BITS(BITS)) U14_MUX_IMAG_4_1
(
    .in_0(x14_i),
    .in_1(x78_i),
    .in_2(x46_i),
    .in_3(x110_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_14_i)
);

MUX_4_1 #(.BITS(BITS)) U15_MUX_IMAG_4_1
(
    .in_0(x30_i),
    .in_1(x94_i),
    .in_2(x62_i),
    .in_3(x126_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_15_i)
);

MUX_4_1 #(.BITS(BITS)) U16_MUX_IMAG_4_1
(
    .in_0(x1_i),
    .in_1(x65_i),
    .in_2(x33_i),
    .in_3(x97_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_16_i)
);

MUX_4_1 #(.BITS(BITS)) U17_MUX_IMAG_4_1
(
    .in_0(x17_i),
    .in_1(x81_i),
    .in_2(x49_i),
    .in_3(x113_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_17_i)
);

MUX_4_1 #(.BITS(BITS)) U18_MUX_IMAG_4_1
(
    .in_0(x9_i),
    .in_1(x73_i),
    .in_2(x41_i),
    .in_3(x105_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_18_i)
);

MUX_4_1 #(.BITS(BITS)) U19_MUX_IMAG_4_1
(
    .in_0(x25_i),
    .in_1(x89_i),
    .in_2(x57_i),
    .in_3(x121_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_19_i)
);

MUX_4_1 #(.BITS(BITS)) U20_MUX_IMAG_4_1
(
    .in_0(x5_i),
    .in_1(x69_i),
    .in_2(x37_i),
    .in_3(x101_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_20_i)
);

MUX_4_1 #(.BITS(BITS)) U21_MUX_IMAG_4_1
(
    .in_0(x21_i),
    .in_1(x85_i),
    .in_2(x53_i),
    .in_3(x117_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_21_i)
);

MUX_4_1 #(.BITS(BITS)) U22_MUX_IMAG_4_1
(
    .in_0(x13_i),
    .in_1(x77_i),
    .in_2(x45_i),
    .in_3(x109_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_22_i)
);

MUX_4_1 #(.BITS(BITS)) U23_MUX_IMAG_4_1
(
    .in_0(x29_i),
    .in_1(x93_i),
    .in_2(x61_i),
    .in_3(x125_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_23_i)
);

MUX_4_1 #(.BITS(BITS)) U24_MUX_IMAG_4_1
(
    .in_0(x3_i),
    .in_1(x67_i),
    .in_2(x35_i),
    .in_3(x99_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_24_i)
);

MUX_4_1 #(.BITS(BITS)) U25_MUX_IMAG_4_1
(
    .in_0(x19_i),
    .in_1(x83_i),
    .in_2(x51_i),
    .in_3(x115_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_25_i)
);

MUX_4_1 #(.BITS(BITS)) U26_MUX_IMAG_4_1
(
    .in_0(x11_i),
    .in_1(x75_i),
    .in_2(x43_i),
    .in_3(x107_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_26_i)
);

MUX_4_1 #(.BITS(BITS)) U27_MUX_IMAG_4_1
(
    .in_0(x27_i),
    .in_1(x91_i),
    .in_2(x59_i),
    .in_3(x123_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_27_i)
);

MUX_4_1 #(.BITS(BITS)) U28_MUX_IMAG_4_1
(
    .in_0(x7_i),
    .in_1(x71_i),
    .in_2(x39_i),
    .in_3(x103_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_28_i)
);

MUX_4_1 #(.BITS(BITS)) U29_MUX_IMAG_4_1
(
    .in_0(x23_i),
    .in_1(x87_i),
    .in_2(x55_i),
    .in_3(x119_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_29_i)
);

MUX_4_1 #(.BITS(BITS)) U30_MUX_IMAG_4_1
(
    .in_0(x15_i),
    .in_1(x79_i),
    .in_2(x47_i),
    .in_3(x111_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_30_i)
);

MUX_4_1 #(.BITS(BITS)) U31_MUX_IMAG_4_1
(
    .in_0(x31_i),
    .in_1(x95_i),
    .in_2(x63_i),
    .in_3(x127_i),
    .selection_line(sel_output_4x1),
    .out(mux4_mux2_31_i)
);







assign X0_r = U0_REAL_MEMORY.locations[0] ;
assign X64_r = U0_REAL_MEMORY.locations[1] ;
assign X1_r = U0_REAL_MEMORY.locations[2] ;
assign X65_r = U0_REAL_MEMORY.locations[3] ;
assign X2_r = U1_REAL_MEMORY.locations[0] ;
assign X66_r = U1_REAL_MEMORY.locations[1] ;
assign X3_r = U1_REAL_MEMORY.locations[2] ;
assign X67_r = U1_REAL_MEMORY.locations[3] ;
assign X4_r = U2_REAL_MEMORY.locations[0] ;
assign X68_r = U2_REAL_MEMORY.locations[1] ;
assign X5_r = U2_REAL_MEMORY.locations[2] ;
assign X69_r = U2_REAL_MEMORY.locations[3] ;
assign X6_r = U3_REAL_MEMORY.locations[0] ;
assign X70_r = U3_REAL_MEMORY.locations[1] ;
assign X7_r = U3_REAL_MEMORY.locations[2] ;
assign X71_r = U3_REAL_MEMORY.locations[3] ;
assign X8_r = U4_REAL_MEMORY.locations[0] ;
assign X72_r = U4_REAL_MEMORY.locations[1] ;
assign X9_r = U4_REAL_MEMORY.locations[2] ;
assign X73_r = U4_REAL_MEMORY.locations[3] ;
assign X10_r = U5_REAL_MEMORY.locations[0] ;
assign X74_r = U5_REAL_MEMORY.locations[1] ;
assign X11_r = U5_REAL_MEMORY.locations[2] ;
assign X75_r = U5_REAL_MEMORY.locations[3] ;
assign X12_r = U6_REAL_MEMORY.locations[0] ;
assign X76_r = U6_REAL_MEMORY.locations[1] ;
assign X13_r = U6_REAL_MEMORY.locations[2] ;
assign X77_r = U6_REAL_MEMORY.locations[3] ;
assign X14_r = U7_REAL_MEMORY.locations[0] ;
assign X78_r = U7_REAL_MEMORY.locations[1] ;
assign X15_r = U7_REAL_MEMORY.locations[2] ;
assign X79_r = U7_REAL_MEMORY.locations[3] ;
assign X16_r = U8_REAL_MEMORY.locations[0] ;
assign X80_r = U8_REAL_MEMORY.locations[1] ;
assign X17_r = U8_REAL_MEMORY.locations[2] ;
assign X81_r = U8_REAL_MEMORY.locations[3] ;
assign X18_r = U9_REAL_MEMORY.locations[0] ;
assign X82_r = U9_REAL_MEMORY.locations[1] ;
assign X19_r = U9_REAL_MEMORY.locations[2] ;
assign X83_r = U9_REAL_MEMORY.locations[3] ;
assign X20_r = U10_REAL_MEMORY.locations[0] ;
assign X84_r = U10_REAL_MEMORY.locations[1] ;
assign X21_r = U10_REAL_MEMORY.locations[2] ;
assign X85_r = U10_REAL_MEMORY.locations[3] ;
assign X22_r = U11_REAL_MEMORY.locations[0] ;
assign X86_r = U11_REAL_MEMORY.locations[1] ;
assign X23_r = U11_REAL_MEMORY.locations[2] ;
assign X87_r = U11_REAL_MEMORY.locations[3] ;
assign X24_r = U12_REAL_MEMORY.locations[0] ;
assign X88_r = U12_REAL_MEMORY.locations[1] ;
assign X25_r = U12_REAL_MEMORY.locations[2] ;
assign X89_r = U12_REAL_MEMORY.locations[3] ;
assign X26_r = U13_REAL_MEMORY.locations[0] ;
assign X90_r = U13_REAL_MEMORY.locations[1] ;
assign X27_r = U13_REAL_MEMORY.locations[2] ;
assign X91_r = U13_REAL_MEMORY.locations[3] ;
assign X28_r = U14_REAL_MEMORY.locations[0] ;
assign X92_r = U14_REAL_MEMORY.locations[1] ;
assign X29_r = U14_REAL_MEMORY.locations[2] ;
assign X93_r = U14_REAL_MEMORY.locations[3] ;
assign X30_r = U15_REAL_MEMORY.locations[0] ;
assign X94_r = U15_REAL_MEMORY.locations[1] ;
assign X31_r = U15_REAL_MEMORY.locations[2] ;
assign X95_r = U15_REAL_MEMORY.locations[3] ;
assign X32_r = U16_REAL_MEMORY.locations[0] ;
assign X96_r = U16_REAL_MEMORY.locations[1] ;
assign X33_r = U16_REAL_MEMORY.locations[2] ;
assign X97_r = U16_REAL_MEMORY.locations[3] ;
assign X34_r = U17_REAL_MEMORY.locations[0] ;
assign X98_r = U17_REAL_MEMORY.locations[1] ;
assign X35_r = U17_REAL_MEMORY.locations[2] ;
assign X99_r = U17_REAL_MEMORY.locations[3] ;
assign X36_r = U18_REAL_MEMORY.locations[0] ;
assign X100_r = U18_REAL_MEMORY.locations[1] ;
assign X37_r = U18_REAL_MEMORY.locations[2] ;
assign X101_r = U18_REAL_MEMORY.locations[3] ;
assign X38_r = U19_REAL_MEMORY.locations[0] ;
assign X102_r = U19_REAL_MEMORY.locations[1] ;
assign X39_r = U19_REAL_MEMORY.locations[2] ;
assign X103_r = U19_REAL_MEMORY.locations[3] ;
assign X40_r = U20_REAL_MEMORY.locations[0] ;
assign X104_r = U20_REAL_MEMORY.locations[1] ;
assign X41_r = U20_REAL_MEMORY.locations[2] ;
assign X105_r = U20_REAL_MEMORY.locations[3] ;
assign X42_r = U21_REAL_MEMORY.locations[0] ;
assign X106_r = U21_REAL_MEMORY.locations[1] ;
assign X43_r = U21_REAL_MEMORY.locations[2] ;
assign X107_r = U21_REAL_MEMORY.locations[3] ;
assign X44_r = U22_REAL_MEMORY.locations[0] ;
assign X108_r = U22_REAL_MEMORY.locations[1] ;
assign X45_r = U22_REAL_MEMORY.locations[2] ;
assign X109_r = U22_REAL_MEMORY.locations[3] ;
assign X46_r = U23_REAL_MEMORY.locations[0] ;
assign X110_r = U23_REAL_MEMORY.locations[1] ;
assign X47_r = U23_REAL_MEMORY.locations[2] ;
assign X111_r = U23_REAL_MEMORY.locations[3] ;
assign X48_r = U24_REAL_MEMORY.locations[0] ;
assign X112_r = U24_REAL_MEMORY.locations[1] ;
assign X49_r = U24_REAL_MEMORY.locations[2] ;
assign X113_r = U24_REAL_MEMORY.locations[3] ;
assign X50_r = U25_REAL_MEMORY.locations[0] ;
assign X114_r = U25_REAL_MEMORY.locations[1] ;
assign X51_r = U25_REAL_MEMORY.locations[2] ;
assign X115_r = U25_REAL_MEMORY.locations[3] ;
assign X52_r = U26_REAL_MEMORY.locations[0] ;
assign X116_r = U26_REAL_MEMORY.locations[1] ;
assign X53_r = U26_REAL_MEMORY.locations[2] ;
assign X117_r = U26_REAL_MEMORY.locations[3] ;
assign X54_r = U27_REAL_MEMORY.locations[0] ;
assign X118_r = U27_REAL_MEMORY.locations[1] ;
assign X55_r = U27_REAL_MEMORY.locations[2] ;
assign X119_r = U27_REAL_MEMORY.locations[3] ;
assign X56_r = U28_REAL_MEMORY.locations[0] ;
assign X120_r = U28_REAL_MEMORY.locations[1] ;
assign X57_r = U28_REAL_MEMORY.locations[2] ;
assign X121_r = U28_REAL_MEMORY.locations[3] ;
assign X58_r = U29_REAL_MEMORY.locations[0] ;
assign X122_r = U29_REAL_MEMORY.locations[1] ;
assign X59_r = U29_REAL_MEMORY.locations[2] ;
assign X123_r = U29_REAL_MEMORY.locations[3] ;
assign X60_r = U30_REAL_MEMORY.locations[0] ;
assign X124_r = U30_REAL_MEMORY.locations[1] ;
assign X61_r = U30_REAL_MEMORY.locations[2] ;
assign X125_r = U30_REAL_MEMORY.locations[3] ;
assign X62_r = U31_REAL_MEMORY.locations[0] ;
assign X126_r = U31_REAL_MEMORY.locations[1] ;
assign X63_r = U31_REAL_MEMORY.locations[2] ;
assign X127_r = U31_REAL_MEMORY.locations[3] ;

assign X0_i = U0_IMAG_MEMORY.locations[0] ;
assign X64_i = U0_IMAG_MEMORY.locations[1] ;
assign X1_i = U0_IMAG_MEMORY.locations[2] ;
assign X65_i = U0_IMAG_MEMORY.locations[3] ;
assign X2_i = U1_IMAG_MEMORY.locations[0] ;
assign X66_i = U1_IMAG_MEMORY.locations[1] ;
assign X3_i = U1_IMAG_MEMORY.locations[2] ;
assign X67_i = U1_IMAG_MEMORY.locations[3] ;
assign X4_i = U2_IMAG_MEMORY.locations[0] ;
assign X68_i = U2_IMAG_MEMORY.locations[1] ;
assign X5_i = U2_IMAG_MEMORY.locations[2] ;
assign X69_i = U2_IMAG_MEMORY.locations[3] ;
assign X6_i = U3_IMAG_MEMORY.locations[0] ;
assign X70_i = U3_IMAG_MEMORY.locations[1] ;
assign X7_i = U3_IMAG_MEMORY.locations[2] ;
assign X71_i = U3_IMAG_MEMORY.locations[3] ;
assign X8_i = U4_IMAG_MEMORY.locations[0] ;
assign X72_i = U4_IMAG_MEMORY.locations[1] ;
assign X9_i = U4_IMAG_MEMORY.locations[2] ;
assign X73_i = U4_IMAG_MEMORY.locations[3] ;
assign X10_i = U5_IMAG_MEMORY.locations[0] ;
assign X74_i = U5_IMAG_MEMORY.locations[1] ;
assign X11_i = U5_IMAG_MEMORY.locations[2] ;
assign X75_i = U5_IMAG_MEMORY.locations[3] ;
assign X12_i = U6_IMAG_MEMORY.locations[0] ;
assign X76_i = U6_IMAG_MEMORY.locations[1] ;
assign X13_i = U6_IMAG_MEMORY.locations[2] ;
assign X77_i = U6_IMAG_MEMORY.locations[3] ;
assign X14_i = U7_IMAG_MEMORY.locations[0] ;
assign X78_i = U7_IMAG_MEMORY.locations[1] ;
assign X15_i = U7_IMAG_MEMORY.locations[2] ;
assign X79_i = U7_IMAG_MEMORY.locations[3] ;
assign X16_i = U8_IMAG_MEMORY.locations[0] ;
assign X80_i = U8_IMAG_MEMORY.locations[1] ;
assign X17_i = U8_IMAG_MEMORY.locations[2] ;
assign X81_i = U8_IMAG_MEMORY.locations[3] ;
assign X18_i = U9_IMAG_MEMORY.locations[0] ;
assign X82_i = U9_IMAG_MEMORY.locations[1] ;
assign X19_i = U9_IMAG_MEMORY.locations[2] ;
assign X83_i = U9_IMAG_MEMORY.locations[3] ;
assign X20_i = U10_IMAG_MEMORY.locations[0] ;
assign X84_i = U10_IMAG_MEMORY.locations[1] ;
assign X21_i = U10_IMAG_MEMORY.locations[2] ;
assign X85_i = U10_IMAG_MEMORY.locations[3] ;
assign X22_i = U11_IMAG_MEMORY.locations[0] ;
assign X86_i = U11_IMAG_MEMORY.locations[1] ;
assign X23_i = U11_IMAG_MEMORY.locations[2] ;
assign X87_i = U11_IMAG_MEMORY.locations[3] ;
assign X24_i = U12_IMAG_MEMORY.locations[0] ;
assign X88_i = U12_IMAG_MEMORY.locations[1] ;
assign X25_i = U12_IMAG_MEMORY.locations[2] ;
assign X89_i = U12_IMAG_MEMORY.locations[3] ;
assign X26_i = U13_IMAG_MEMORY.locations[0] ;
assign X90_i = U13_IMAG_MEMORY.locations[1] ;
assign X27_i = U13_IMAG_MEMORY.locations[2] ;
assign X91_i = U13_IMAG_MEMORY.locations[3] ;
assign X28_i = U14_IMAG_MEMORY.locations[0] ;
assign X92_i = U14_IMAG_MEMORY.locations[1] ;
assign X29_i = U14_IMAG_MEMORY.locations[2] ;
assign X93_i = U14_IMAG_MEMORY.locations[3] ;
assign X30_i = U15_IMAG_MEMORY.locations[0] ;
assign X94_i = U15_IMAG_MEMORY.locations[1] ;
assign X31_i = U15_IMAG_MEMORY.locations[2] ;
assign X95_i = U15_IMAG_MEMORY.locations[3] ;
assign X32_i = U16_IMAG_MEMORY.locations[0] ;
assign X96_i = U16_IMAG_MEMORY.locations[1] ;
assign X33_i = U16_IMAG_MEMORY.locations[2] ;
assign X97_i = U16_IMAG_MEMORY.locations[3] ;
assign X34_i = U17_IMAG_MEMORY.locations[0] ;
assign X98_i = U17_IMAG_MEMORY.locations[1] ;
assign X35_i = U17_IMAG_MEMORY.locations[2] ;
assign X99_i = U17_IMAG_MEMORY.locations[3] ;
assign X36_i = U18_IMAG_MEMORY.locations[0] ;
assign X100_i = U18_IMAG_MEMORY.locations[1] ;
assign X37_i = U18_IMAG_MEMORY.locations[2] ;
assign X101_i = U18_IMAG_MEMORY.locations[3] ;
assign X38_i = U19_IMAG_MEMORY.locations[0] ;
assign X102_i = U19_IMAG_MEMORY.locations[1] ;
assign X39_i = U19_IMAG_MEMORY.locations[2] ;
assign X103_i = U19_IMAG_MEMORY.locations[3] ;
assign X40_i = U20_IMAG_MEMORY.locations[0] ;
assign X104_i = U20_IMAG_MEMORY.locations[1] ;
assign X41_i = U20_IMAG_MEMORY.locations[2] ;
assign X105_i = U20_IMAG_MEMORY.locations[3] ;
assign X42_i = U21_IMAG_MEMORY.locations[0] ;
assign X106_i = U21_IMAG_MEMORY.locations[1] ;
assign X43_i = U21_IMAG_MEMORY.locations[2] ;
assign X107_i = U21_IMAG_MEMORY.locations[3] ;
assign X44_i = U22_IMAG_MEMORY.locations[0] ;
assign X108_i = U22_IMAG_MEMORY.locations[1] ;
assign X45_i = U22_IMAG_MEMORY.locations[2] ;
assign X109_i = U22_IMAG_MEMORY.locations[3] ;
assign X46_i = U23_IMAG_MEMORY.locations[0] ;
assign X110_i = U23_IMAG_MEMORY.locations[1] ;
assign X47_i = U23_IMAG_MEMORY.locations[2] ;
assign X111_i = U23_IMAG_MEMORY.locations[3] ;
assign X48_i = U24_IMAG_MEMORY.locations[0] ;
assign X112_i = U24_IMAG_MEMORY.locations[1] ;
assign X49_i = U24_IMAG_MEMORY.locations[2] ;
assign X113_i = U24_IMAG_MEMORY.locations[3] ;
assign X50_i = U25_IMAG_MEMORY.locations[0] ;
assign X114_i = U25_IMAG_MEMORY.locations[1] ;
assign X51_i = U25_IMAG_MEMORY.locations[2] ;
assign X115_i = U25_IMAG_MEMORY.locations[3] ;
assign X52_i = U26_IMAG_MEMORY.locations[0] ;
assign X116_i = U26_IMAG_MEMORY.locations[1] ;
assign X53_i = U26_IMAG_MEMORY.locations[2] ;
assign X117_i = U26_IMAG_MEMORY.locations[3] ;
assign X54_i = U27_IMAG_MEMORY.locations[0] ;
assign X118_i = U27_IMAG_MEMORY.locations[1] ;
assign X55_i = U27_IMAG_MEMORY.locations[2] ;
assign X119_i = U27_IMAG_MEMORY.locations[3] ;
assign X56_i = U28_IMAG_MEMORY.locations[0] ;
assign X120_i = U28_IMAG_MEMORY.locations[1] ;
assign X57_i = U28_IMAG_MEMORY.locations[2] ;
assign X121_i = U28_IMAG_MEMORY.locations[3] ;
assign X58_i = U29_IMAG_MEMORY.locations[0] ;
assign X122_i = U29_IMAG_MEMORY.locations[1] ;
assign X59_i = U29_IMAG_MEMORY.locations[2] ;
assign X123_i = U29_IMAG_MEMORY.locations[3] ;
assign X60_i = U30_IMAG_MEMORY.locations[0] ;
assign X124_i = U30_IMAG_MEMORY.locations[1] ;
assign X61_i = U30_IMAG_MEMORY.locations[2] ;
assign X125_i = U30_IMAG_MEMORY.locations[3] ;
assign X62_i = U31_IMAG_MEMORY.locations[0] ;
assign X126_i = U31_IMAG_MEMORY.locations[1] ;
assign X63_i = U31_IMAG_MEMORY.locations[2] ;
assign X127_i = U31_IMAG_MEMORY.locations[3] ;


endmodule
