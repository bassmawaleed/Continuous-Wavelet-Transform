
`timescale 1ns/1ps

module cwt_top_module_tb();
	
	
	/* Parameters */
	parameter Clock_Period = 4 ;
	parameter BITS =16;

     integer inputs ;


	/* FIRST : Define the testbench signals */
	///////////// Inputs /////////////
    reg ready_inputs_tb ;
    reg clk_tb;
    reg rst_tb;
    reg [1:0] read_scale_ram_addresses;
    reg [BITS-1 : 0 ] x0_r_tb ;
    reg [BITS-1 : 0 ] x0_i_tb ;
    reg [BITS-1 : 0 ] x1_r_tb ;
    reg [BITS-1 : 0 ] x1_i_tb ;
    reg [BITS-1 : 0 ] x2_r_tb ;
    reg [BITS-1 : 0 ] x2_i_tb;
    reg [BITS-1 : 0 ] x3_r_tb ;
    reg [BITS-1 : 0 ] x3_i_tb ;
    reg [BITS-1 : 0 ] x4_r_tb ;
    reg [BITS-1 : 0 ] x4_i_tb ;
    reg [BITS-1 : 0 ] x5_r_tb ;
    reg [BITS-1 : 0 ] x5_i_tb ;
    reg [BITS-1 : 0 ] x6_r_tb ;
    reg [BITS-1 : 0 ] x6_i_tb ;
    reg[BITS-1 : 0 ] x7_r_tb ;
    reg [BITS-1 : 0 ] x7_i_tb;
    reg [BITS-1 : 0 ] x8_r_tb;
    reg [BITS-1 : 0 ] x8_i_tb;
    reg [BITS-1 : 0 ] x9_r_tb;
    reg [BITS-1 : 0 ] x9_i_tb;
    reg [BITS-1 : 0 ] x10_r_tb;
    reg [BITS-1 : 0 ] x10_i_tb;
    reg [BITS-1 : 0 ] x11_r_tb;
    reg [BITS-1 : 0 ] x11_i_tb;
    reg [BITS-1 : 0 ] x12_r_tb;
    reg [BITS-1 : 0 ] x12_i_tb;
    reg [BITS-1 : 0 ] x13_r_tb;
    reg [BITS-1 : 0 ] x13_i_tb;
    reg [BITS-1 : 0 ] x14_r_tb;
    reg [BITS-1 : 0 ] x14_i_tb;
    reg [BITS-1 : 0 ] x15_r_tb;
    reg [BITS-1 : 0 ] x15_i_tb;
    reg [BITS-1 : 0 ] x16_r_tb ;
    reg [BITS-1 : 0 ] x16_i_tb ;
    reg [BITS-1 : 0 ] x17_r_tb ;
    reg [BITS-1 : 0 ] x17_i_tb ;
    reg [BITS-1 : 0 ] x18_r_tb ;
    reg [BITS-1 : 0 ] x18_i_tb;
    reg [BITS-1 : 0 ] x19_r_tb ;
    reg [BITS-1 : 0 ] x19_i_tb ;
    reg [BITS-1 : 0 ] x20_r_tb ;
    reg [BITS-1 : 0 ] x20_i_tb ;
    reg [BITS-1 : 0 ] x21_r_tb ;
    reg [BITS-1 : 0 ] x21_i_tb ;
    reg [BITS-1 : 0 ] x22_r_tb ;
    reg [BITS-1 : 0 ] x22_i_tb ;
    reg [BITS-1 : 0 ] x23_r_tb ;
    reg [BITS-1 : 0 ] x23_i_tb ;
    reg[BITS-1 : 0 ] x24_r_tb ;
    reg [BITS-1 : 0 ] x24_i_tb;
    reg [BITS-1 : 0 ] x25_r_tb;
    reg [BITS-1 : 0 ] x25_i_tb;
    reg [BITS-1 : 0 ] x26_r_tb;
    reg [BITS-1 : 0 ] x26_i_tb;
    reg [BITS-1 : 0 ] x27_r_tb;
    reg [BITS-1 : 0 ] x27_i_tb;
    reg [BITS-1 : 0 ] x28_r_tb;
    reg [BITS-1 : 0 ] x28_i_tb;
    reg [BITS-1 : 0 ] x29_r_tb;
    reg [BITS-1 : 0 ] x29_i_tb;
    reg [BITS-1 : 0 ] x30_r_tb;
    reg [BITS-1 : 0 ] x30_i_tb;
    reg [BITS-1 : 0 ] x31_r_tb;
    reg[BITS-1 : 0 ] x31_i_tb;
    reg [BITS-1 : 0 ] x32_r_tb;
    reg [BITS-1 : 0 ] x32_i_tb;
    reg [BITS-1 : 0 ] x33_r_tb ;
    reg [BITS-1 : 0 ] x33_i_tb ;
    reg [BITS-1 : 0 ] x34_r_tb ;
    reg [BITS-1 : 0 ] x34_i_tb ;
    reg [BITS-1 : 0 ] x35_r_tb ;
    reg [BITS-1 : 0 ] x35_i_tb;
    reg [BITS-1 : 0 ] x36_r_tb ;
    reg [BITS-1 : 0 ] x36_i_tb ;
    reg [BITS-1 : 0 ] x37_r_tb ;
    reg [BITS-1 : 0 ] x37_i_tb ;
    reg [BITS-1 : 0 ] x38_r_tb ;
    reg [BITS-1 : 0 ] x38_i_tb ;
    reg [BITS-1 : 0 ] x39_r_tb ;
    reg [BITS-1 : 0 ] x39_i_tb ;
    reg[BITS-1 : 0 ] x40_r_tb ;
    reg [BITS-1 : 0 ] x40_i_tb;
    reg [BITS-1 : 0 ] x41_r_tb;
    reg [BITS-1 : 0 ] x41_i_tb;
    reg [BITS-1 : 0 ] x42_r_tb;
    reg [BITS-1 : 0 ] x42_i_tb;
    reg [BITS-1 : 0 ] x43_r_tb;
    reg [BITS-1 : 0 ] x43_i_tb;
    reg [BITS-1 : 0 ] x44_r_tb;
    reg [BITS-1 : 0 ] x44_i_tb;
    reg [BITS-1 : 0 ] x45_r_tb;
    reg [BITS-1 : 0 ] x45_i_tb;
    reg [BITS-1 : 0 ] x46_r_tb;
    reg [BITS-1 : 0 ] x46_i_tb;
    reg [BITS-1 : 0 ] x47_r_tb;
    reg[BITS-1 : 0 ] x47_i_tb;
    reg [BITS-1 : 0 ] x48_r_tb;
    reg [BITS-1 : 0 ] x48_i_tb;
    reg [BITS-1 : 0 ] x49_r_tb ;
    reg [BITS-1 : 0 ] x49_i_tb ;
    reg [BITS-1 : 0 ] x50_r_tb ;
    reg [BITS-1 : 0 ] x50_i_tb ;
    reg [BITS-1 : 0 ] x51_r_tb ;
    reg [BITS-1 : 0 ] x51_i_tb;
    reg [BITS-1 : 0 ] x52_r_tb ;
    reg [BITS-1 : 0 ] x52_i_tb ;
    reg [BITS-1 : 0 ] x53_r_tb ;
    reg [BITS-1 : 0 ] x53_i_tb ;
    reg [BITS-1 : 0 ] x54_r_tb ;
    reg [BITS-1 : 0 ] x54_i_tb ;
    reg [BITS-1 : 0 ] x55_r_tb ;
    reg [BITS-1 : 0 ] x55_i_tb ;
    reg[BITS-1 : 0 ] x56_r_tb ;
    reg [BITS-1 : 0 ] x56_i_tb;
    reg [BITS-1 : 0 ] x57_r_tb;
    reg [BITS-1 : 0 ] x57_i_tb;
    reg [BITS-1 : 0 ] x58_r_tb;
    reg [BITS-1 : 0 ] x58_i_tb;
    reg [BITS-1 : 0 ] x59_r_tb;
    reg [BITS-1 : 0 ] x59_i_tb;
    reg [BITS-1 : 0 ] x60_r_tb;
    reg [BITS-1 : 0 ] x60_i_tb;
    reg [BITS-1 : 0 ] x61_r_tb;
    reg [BITS-1 : 0 ] x61_i_tb;
    reg [BITS-1 : 0 ] x62_r_tb;
    reg [BITS-1 : 0 ] x62_i_tb;
    reg [BITS-1 : 0 ] x63_r_tb;
    reg [BITS-1 : 0 ] x63_i_tb;
    reg [BITS-1 : 0 ] x64_r_tb;
    reg [BITS-1 : 0 ] x64_i_tb;
    reg [BITS-1 : 0 ] x65_r_tb ;
    reg [BITS-1 : 0 ] x65_i_tb ;
    reg [BITS-1 : 0 ] x66_r_tb ;
    reg [BITS-1 : 0 ] x66_i_tb ;
    reg [BITS-1 : 0 ] x67_r_tb ;
    reg [BITS-1 : 0 ] x67_i_tb;
    reg [BITS-1 : 0 ] x68_r_tb ;
    reg  [BITS-1 : 0 ] x68_i_tb ;
    reg [BITS-1 : 0 ] x69_r_tb ;
    reg [BITS-1 : 0 ] x69_i_tb ;
    reg [BITS-1 : 0 ] x70_r_tb ;
    reg [BITS-1 : 0 ] x70_i_tb ;
    reg [BITS-1 : 0 ] x71_r_tb ;
    reg [BITS-1 : 0 ] x71_i_tb ;
    reg [BITS-1 : 0 ] x72_r_tb ;
    reg [BITS-1 : 0 ] x72_i_tb;
    reg [BITS-1 : 0 ] x73_r_tb;
    reg [BITS-1 : 0 ] x73_i_tb;
    reg [BITS-1 : 0 ] x74_r_tb;
    reg [BITS-1 : 0 ] x74_i_tb;
    reg [BITS-1 : 0 ] x75_r_tb;
    reg [BITS-1 : 0 ] x75_i_tb;
    reg [BITS-1 : 0 ] x76_r_tb;
    reg [BITS-1 : 0 ] x76_i_tb;
    reg [BITS-1 : 0 ] x77_r_tb;
    reg [BITS-1 : 0 ] x77_i_tb;
    reg [BITS-1 : 0 ] x78_r_tb;
    reg [BITS-1 : 0 ] x78_i_tb;
    reg [BITS-1 : 0 ] x79_r_tb;
    reg [BITS-1 : 0 ] x79_i_tb;
    reg [BITS-1 : 0 ] x80_r_tb;
    reg [BITS-1 : 0 ] x80_i_tb;
    reg [BITS-1 : 0 ] x81_r_tb ;
    reg [BITS-1 : 0 ] x81_i_tb ;
    reg [BITS-1 : 0 ] x82_r_tb ;
    reg [BITS-1 : 0 ] x82_i_tb ;
    reg [BITS-1 : 0 ] x83_r_tb ;
    reg [BITS-1 : 0 ] x83_i_tb;
    reg [BITS-1 : 0 ] x84_r_tb ;
    reg [BITS-1 : 0 ] x84_i_tb ;
    reg [BITS-1 : 0 ] x85_r_tb ;
    reg [BITS-1 : 0 ] x85_i_tb ;
    reg [BITS-1 : 0 ] x86_r_tb ;
    reg [BITS-1 : 0 ] x86_i_tb ;
    reg [BITS-1 : 0 ] x87_r_tb ;
    reg [BITS-1 : 0 ] x87_i_tb ;
    reg[BITS-1 : 0 ] x88_r_tb ;
    reg [BITS-1 : 0 ] x88_i_tb;
    reg [BITS-1 : 0 ] x89_r_tb;
    reg [BITS-1 : 0 ] x89_i_tb;
    reg [BITS-1 : 0 ] x90_r_tb;
    reg [BITS-1 : 0 ] x90_i_tb;
    reg [BITS-1 : 0 ] x91_r_tb;
    reg [BITS-1 : 0 ] x91_i_tb;
    reg [BITS-1 : 0 ] x92_r_tb;
    reg [BITS-1 : 0 ] x92_i_tb;
    reg [BITS-1 : 0 ] x93_r_tb;
    reg [BITS-1 : 0 ] x93_i_tb;
    reg [BITS-1 : 0 ] x94_r_tb;
    reg [BITS-1 : 0 ] x94_i_tb;
    reg [BITS-1 : 0 ] x95_r_tb;
    reg [BITS-1 : 0 ] x95_i_tb;
    reg [BITS-1 : 0 ] x96_r_tb;
    reg [BITS-1 : 0 ] x96_i_tb;
    reg [BITS-1 : 0 ] x97_r_tb ;
    reg [BITS-1 : 0 ] x97_i_tb ;
    reg [BITS-1 : 0 ] x98_r_tb ;
    reg [BITS-1 : 0 ] x98_i_tb ;
    reg [BITS-1 : 0 ] x99_r_tb ;
    reg [BITS-1 : 0 ] x99_i_tb;
    reg [BITS-1 : 0 ] x100_r_tb ;
    reg [BITS-1 : 0 ] x100_i_tb ;
    reg [BITS-1 : 0 ] x101_r_tb ;
    reg [BITS-1 : 0 ] x101_i_tb ;
    reg [BITS-1 : 0 ] x102_r_tb ;
    reg [BITS-1 : 0 ] x102_i_tb ;
    reg [BITS-1 : 0 ] x103_r_tb ;
    reg [BITS-1 : 0 ] x103_i_tb ;
    reg [BITS-1 : 0 ] x104_r_tb ;
    reg [BITS-1 : 0 ] x104_i_tb;
    reg [BITS-1 : 0 ] x105_r_tb;
    reg [BITS-1 : 0 ] x105_i_tb;
    reg [BITS-1 : 0 ] x106_r_tb;
    reg [BITS-1 : 0 ] x106_i_tb;
    reg [BITS-1 : 0 ] x107_r_tb;
    reg [BITS-1 : 0 ] x107_i_tb;
    reg [BITS-1 : 0 ] x108_r_tb;
    reg [BITS-1 : 0 ] x108_i_tb;
    reg [BITS-1 : 0 ] x109_r_tb;
    reg [BITS-1 : 0 ] x109_i_tb;
    reg [BITS-1 : 0 ] x110_r_tb;
    reg [BITS-1 : 0 ] x110_i_tb;
    reg [BITS-1 : 0 ] x111_r_tb;
    reg [BITS-1 : 0 ] x111_i_tb;
    reg [BITS-1 : 0 ] x112_r_tb;
    reg [BITS-1 : 0 ] x112_i_tb;
    reg [BITS-1 : 0 ] x113_r_tb ;
    reg [BITS-1 : 0 ] x113_i_tb ;
    reg [BITS-1 : 0 ] x114_r_tb ;
    reg [BITS-1 : 0 ] x114_i_tb ;
    reg [BITS-1 : 0 ] x115_r_tb ;
    reg [BITS-1 : 0 ] x115_i_tb;
    reg [BITS-1 : 0 ] x116_r_tb ;
    reg [BITS-1 : 0 ] x116_i_tb ;
    reg [BITS-1 : 0 ] x117_r_tb ;
    reg [BITS-1 : 0 ] x117_i_tb ;
    reg [BITS-1 : 0 ] x118_r_tb ;
    reg [BITS-1 : 0 ] x118_i_tb ;
    reg [BITS-1 : 0 ] x119_r_tb ;
    reg [BITS-1 : 0 ] x119_i_tb ;
    reg [BITS-1 : 0 ] x120_r_tb ;
    reg [BITS-1 : 0 ] x120_i_tb;
    reg [BITS-1 : 0 ] x121_r_tb;
    reg [BITS-1 : 0 ] x121_i_tb;
    reg [BITS-1 : 0 ] x122_r_tb;
    reg [BITS-1 : 0 ] x122_i_tb;
    reg [BITS-1 : 0 ] x123_r_tb;
    reg [BITS-1 : 0 ] x123_i_tb;
    reg [BITS-1 : 0 ] x124_r_tb;
    reg [BITS-1 : 0 ] x124_i_tb;
    reg [BITS-1 : 0 ] x125_r_tb;
    reg [BITS-1 : 0 ] x125_i_tb;
    reg [BITS-1 : 0 ] x126_r_tb;
    reg [BITS-1 : 0 ] x126_i_tb;
    reg [BITS-1 : 0 ] x127_r_tb;
    reg [BITS-1 : 0 ] x127_i_tb;



    wire [BITS-1:0] memory_0_scale_1_real_tb;
    wire [BITS-1:0] memory_1_scale_1_real_tb;
    wire [BITS-1:0] memory_2_scale_1_real_tb;
    wire [BITS-1:0] memory_3_scale_1_real_tb;
    wire [BITS-1:0] memory_4_scale_1_real_tb;
    wire [BITS-1:0] memory_5_scale_1_real_tb;
    wire [BITS-1:0] memory_6_scale_1_real_tb;
    wire [BITS-1:0] memory_7_scale_1_real_tb;
    wire [BITS-1:0] memory_8_scale_1_real_tb;
    wire [BITS-1:0] memory_9_scale_1_real_tb;
    wire [BITS-1:0] memory_10_scale_1_real_tb;
    wire [BITS-1:0] memory_11_scale_1_real_tb;
    wire [BITS-1:0] memory_12_scale_1_real_tb;
    wire [BITS-1:0] memory_13_scale_1_real_tb;
    wire [BITS-1:0] memory_14_scale_1_real_tb;
    wire [BITS-1:0] memory_15_scale_1_real_tb;
    wire [BITS-1:0] memory_16_scale_1_real_tb;
    wire [BITS-1:0] memory_17_scale_1_real_tb;
    wire [BITS-1:0] memory_18_scale_1_real_tb;
    wire [BITS-1:0] memory_19_scale_1_real_tb;
    wire [BITS-1:0] memory_20_scale_1_real_tb;
    wire [BITS-1:0] memory_21_scale_1_real_tb;
    wire [BITS-1:0] memory_22_scale_1_real_tb;
    wire [BITS-1:0] memory_23_scale_1_real_tb;
    wire [BITS-1:0] memory_24_scale_1_real_tb;
    wire [BITS-1:0] memory_25_scale_1_real_tb;
    wire [BITS-1:0] memory_26_scale_1_real_tb;
    wire [BITS-1:0] memory_27_scale_1_real_tb;
    wire [BITS-1:0] memory_28_scale_1_real_tb;
    wire [BITS-1:0] memory_29_scale_1_real_tb;
    wire [BITS-1:0] memory_30_scale_1_real_tb;
    wire [BITS-1:0] memory_31_scale_1_real_tb;
    wire [BITS-1:0] memory_0_scale_2_real_tb;
    wire [BITS-1:0] memory_1_scale_2_real_tb;
    wire [BITS-1:0] memory_2_scale_2_real_tb;
    wire [BITS-1:0] memory_3_scale_2_real_tb;
    wire [BITS-1:0] memory_4_scale_2_real_tb;
    wire [BITS-1:0] memory_5_scale_2_real_tb;
    wire [BITS-1:0] memory_6_scale_2_real_tb;
    wire [BITS-1:0] memory_7_scale_2_real_tb;
    wire [BITS-1:0] memory_8_scale_2_real_tb;
    wire [BITS-1:0] memory_9_scale_2_real_tb;
    wire [BITS-1:0] memory_10_scale_2_real_tb;
    wire [BITS-1:0] memory_11_scale_2_real_tb;
    wire [BITS-1:0] memory_12_scale_2_real_tb;
    wire [BITS-1:0] memory_13_scale_2_real_tb;
    wire [BITS-1:0] memory_14_scale_2_real_tb;
    wire [BITS-1:0] memory_15_scale_2_real_tb;
    wire [BITS-1:0] memory_16_scale_2_real_tb;
    wire [BITS-1:0] memory_17_scale_2_real_tb;
    wire [BITS-1:0] memory_18_scale_2_real_tb;
    wire [BITS-1:0] memory_19_scale_2_real_tb;
    wire [BITS-1:0] memory_20_scale_2_real_tb;
    wire [BITS-1:0] memory_21_scale_2_real_tb;
    wire [BITS-1:0] memory_22_scale_2_real_tb;
    wire [BITS-1:0] memory_23_scale_2_real_tb;
    wire [BITS-1:0] memory_24_scale_2_real_tb;
    wire [BITS-1:0] memory_25_scale_2_real_tb;
    wire [BITS-1:0] memory_26_scale_2_real_tb;
    wire [BITS-1:0] memory_27_scale_2_real_tb;
    wire [BITS-1:0] memory_28_scale_2_real_tb;
    wire [BITS-1:0] memory_29_scale_2_real_tb;
    wire [BITS-1:0] memory_30_scale_2_real_tb;
    wire [BITS-1:0] memory_31_scale_2_real_tb;
    wire [BITS-1:0] memory_0_scale_3_real_tb;
    wire [BITS-1:0] memory_1_scale_3_real_tb;
    wire [BITS-1:0] memory_2_scale_3_real_tb;
    wire [BITS-1:0] memory_3_scale_3_real_tb;
    wire [BITS-1:0] memory_4_scale_3_real_tb;
    wire [BITS-1:0] memory_5_scale_3_real_tb;
    wire [BITS-1:0] memory_6_scale_3_real_tb;
    wire [BITS-1:0] memory_7_scale_3_real_tb;
    wire [BITS-1:0] memory_8_scale_3_real_tb;
    wire [BITS-1:0] memory_9_scale_3_real_tb;
    wire [BITS-1:0] memory_10_scale_3_real_tb;
    wire [BITS-1:0] memory_11_scale_3_real_tb;
    wire [BITS-1:0] memory_12_scale_3_real_tb;
    wire [BITS-1:0] memory_13_scale_3_real_tb;
    wire [BITS-1:0] memory_14_scale_3_real_tb;
    wire [BITS-1:0] memory_15_scale_3_real_tb;
    wire [BITS-1:0] memory_16_scale_3_real_tb;
    wire [BITS-1:0] memory_17_scale_3_real_tb;
    wire [BITS-1:0] memory_18_scale_3_real_tb;
    wire [BITS-1:0] memory_19_scale_3_real_tb;
    wire [BITS-1:0] memory_20_scale_3_real_tb;
    wire [BITS-1:0] memory_21_scale_3_real_tb;
    wire [BITS-1:0] memory_22_scale_3_real_tb;
    wire [BITS-1:0] memory_23_scale_3_real_tb;
    wire [BITS-1:0] memory_24_scale_3_real_tb;
    wire [BITS-1:0] memory_25_scale_3_real_tb;
    wire [BITS-1:0] memory_26_scale_3_real_tb;
    wire [BITS-1:0] memory_27_scale_3_real_tb;
    wire [BITS-1:0] memory_28_scale_3_real_tb;
    wire [BITS-1:0] memory_29_scale_3_real_tb;
    wire [BITS-1:0] memory_30_scale_3_real_tb;
    wire [BITS-1:0] memory_31_scale_3_real_tb;
    wire [BITS-1:0] memory_0_scale_4_real_tb;
    wire [BITS-1:0] memory_1_scale_4_real_tb;
    wire [BITS-1:0] memory_2_scale_4_real_tb;
    wire [BITS-1:0] memory_3_scale_4_real_tb;
    wire [BITS-1:0] memory_4_scale_4_real_tb;
    wire [BITS-1:0] memory_5_scale_4_real_tb;
    wire [BITS-1:0] memory_6_scale_4_real_tb;
    wire [BITS-1:0] memory_7_scale_4_real_tb;
    wire [BITS-1:0] memory_8_scale_4_real_tb;
    wire [BITS-1:0] memory_9_scale_4_real_tb;
    wire [BITS-1:0] memory_10_scale_4_real_tb;
    wire [BITS-1:0] memory_11_scale_4_real_tb;
    wire [BITS-1:0] memory_12_scale_4_real_tb;
    wire [BITS-1:0] memory_13_scale_4_real_tb;
    wire [BITS-1:0] memory_14_scale_4_real_tb;
    wire [BITS-1:0] memory_15_scale_4_real_tb;
    wire [BITS-1:0] memory_16_scale_4_real_tb;
    wire [BITS-1:0] memory_17_scale_4_real_tb;
    wire [BITS-1:0] memory_18_scale_4_real_tb;
    wire [BITS-1:0] memory_19_scale_4_real_tb;
    wire [BITS-1:0] memory_20_scale_4_real_tb;
    wire [BITS-1:0] memory_21_scale_4_real_tb;
    wire [BITS-1:0] memory_22_scale_4_real_tb;
    wire [BITS-1:0] memory_23_scale_4_real_tb;
    wire [BITS-1:0] memory_24_scale_4_real_tb;
    wire [BITS-1:0] memory_25_scale_4_real_tb;
    wire [BITS-1:0] memory_26_scale_4_real_tb;
    wire [BITS-1:0] memory_27_scale_4_real_tb;
    wire [BITS-1:0] memory_28_scale_4_real_tb;
    wire [BITS-1:0] memory_29_scale_4_real_tb;
    wire [BITS-1:0] memory_30_scale_4_real_tb;
    wire [BITS-1:0] memory_31_scale_4_real_tb;
    wire [BITS-1:0] memory_0_scale_5_real_tb;
    wire [BITS-1:0] memory_1_scale_5_real_tb;
    wire [BITS-1:0] memory_2_scale_5_real_tb;
    wire [BITS-1:0] memory_3_scale_5_real_tb;
    wire [BITS-1:0] memory_4_scale_5_real_tb;
    wire [BITS-1:0] memory_5_scale_5_real_tb;
    wire [BITS-1:0] memory_6_scale_5_real_tb;
    wire [BITS-1:0] memory_7_scale_5_real_tb;
    wire [BITS-1:0] memory_8_scale_5_real_tb;
    wire [BITS-1:0] memory_9_scale_5_real_tb;
    wire [BITS-1:0] memory_10_scale_5_real_tb;
    wire [BITS-1:0] memory_11_scale_5_real_tb;
    wire [BITS-1:0] memory_12_scale_5_real_tb;
    wire [BITS-1:0] memory_13_scale_5_real_tb;
    wire [BITS-1:0] memory_14_scale_5_real_tb;
    wire [BITS-1:0] memory_15_scale_5_real_tb;
    wire [BITS-1:0] memory_16_scale_5_real_tb;
    wire [BITS-1:0] memory_17_scale_5_real_tb;
    wire [BITS-1:0] memory_18_scale_5_real_tb;
    wire [BITS-1:0] memory_19_scale_5_real_tb;
    wire [BITS-1:0] memory_20_scale_5_real_tb;
    wire [BITS-1:0] memory_21_scale_5_real_tb;
    wire [BITS-1:0] memory_22_scale_5_real_tb;
    wire [BITS-1:0] memory_23_scale_5_real_tb;
    wire [BITS-1:0] memory_24_scale_5_real_tb;
    wire [BITS-1:0] memory_25_scale_5_real_tb;
    wire [BITS-1:0] memory_26_scale_5_real_tb;
    wire [BITS-1:0] memory_27_scale_5_real_tb;
    wire [BITS-1:0] memory_28_scale_5_real_tb;
    wire [BITS-1:0] memory_29_scale_5_real_tb;
    wire [BITS-1:0] memory_30_scale_5_real_tb;
    wire [BITS-1:0] memory_31_scale_5_real_tb;
    wire [BITS-1:0] memory_0_scale_6_real_tb;
    wire [BITS-1:0] memory_1_scale_6_real_tb;
    wire [BITS-1:0] memory_2_scale_6_real_tb;
    wire [BITS-1:0] memory_3_scale_6_real_tb;
    wire [BITS-1:0] memory_4_scale_6_real_tb;
    wire [BITS-1:0] memory_5_scale_6_real_tb;
    wire [BITS-1:0] memory_6_scale_6_real_tb;
    wire [BITS-1:0] memory_7_scale_6_real_tb;
    wire [BITS-1:0] memory_8_scale_6_real_tb;
    wire [BITS-1:0] memory_9_scale_6_real_tb;
    wire [BITS-1:0] memory_10_scale_6_real_tb;
    wire [BITS-1:0] memory_11_scale_6_real_tb;
    wire [BITS-1:0] memory_12_scale_6_real_tb;
    wire [BITS-1:0] memory_13_scale_6_real_tb;
    wire [BITS-1:0] memory_14_scale_6_real_tb;
    wire [BITS-1:0] memory_15_scale_6_real_tb;
    wire [BITS-1:0] memory_16_scale_6_real_tb;
    wire [BITS-1:0] memory_17_scale_6_real_tb;
    wire [BITS-1:0] memory_18_scale_6_real_tb;
    wire [BITS-1:0] memory_19_scale_6_real_tb;
    wire [BITS-1:0] memory_20_scale_6_real_tb;
    wire [BITS-1:0] memory_21_scale_6_real_tb;
    wire [BITS-1:0] memory_22_scale_6_real_tb;
    wire [BITS-1:0] memory_23_scale_6_real_tb;
    wire [BITS-1:0] memory_24_scale_6_real_tb;
    wire [BITS-1:0] memory_25_scale_6_real_tb;
    wire [BITS-1:0] memory_26_scale_6_real_tb;
    wire [BITS-1:0] memory_27_scale_6_real_tb;
    wire [BITS-1:0] memory_28_scale_6_real_tb;
    wire [BITS-1:0] memory_29_scale_6_real_tb;
    wire [BITS-1:0] memory_30_scale_6_real_tb;
    wire [BITS-1:0] memory_31_scale_6_real_tb;
    wire [BITS-1:0] memory_0_scale_7_real_tb;
    wire [BITS-1:0] memory_1_scale_7_real_tb;
    wire [BITS-1:0] memory_2_scale_7_real_tb;
    wire [BITS-1:0] memory_3_scale_7_real_tb;
    wire [BITS-1:0] memory_4_scale_7_real_tb;
    wire [BITS-1:0] memory_5_scale_7_real_tb;
    wire [BITS-1:0] memory_6_scale_7_real_tb;
    wire [BITS-1:0] memory_7_scale_7_real_tb;
    wire [BITS-1:0] memory_8_scale_7_real_tb;
    wire [BITS-1:0] memory_9_scale_7_real_tb;
    wire [BITS-1:0] memory_10_scale_7_real_tb;
    wire [BITS-1:0] memory_11_scale_7_real_tb;
    wire [BITS-1:0] memory_12_scale_7_real_tb;
    wire [BITS-1:0] memory_13_scale_7_real_tb;
    wire [BITS-1:0] memory_14_scale_7_real_tb;
    wire [BITS-1:0] memory_15_scale_7_real_tb;
    wire [BITS-1:0] memory_16_scale_7_real_tb;
    wire [BITS-1:0] memory_17_scale_7_real_tb;
    wire [BITS-1:0] memory_18_scale_7_real_tb;
    wire [BITS-1:0] memory_19_scale_7_real_tb;
    wire [BITS-1:0] memory_20_scale_7_real_tb;
    wire [BITS-1:0] memory_21_scale_7_real_tb;
    wire [BITS-1:0] memory_22_scale_7_real_tb;
    wire [BITS-1:0] memory_23_scale_7_real_tb;
    wire [BITS-1:0] memory_24_scale_7_real_tb;
    wire [BITS-1:0] memory_25_scale_7_real_tb;
    wire [BITS-1:0] memory_26_scale_7_real_tb;
    wire [BITS-1:0] memory_27_scale_7_real_tb;
    wire [BITS-1:0] memory_28_scale_7_real_tb;
    wire [BITS-1:0] memory_29_scale_7_real_tb;
    wire [BITS-1:0] memory_30_scale_7_real_tb;
    wire [BITS-1:0] memory_31_scale_7_real_tb;
    wire [BITS-1:0] memory_0_scale_8_real_tb;
    wire [BITS-1:0] memory_1_scale_8_real_tb;
    wire [BITS-1:0] memory_2_scale_8_real_tb;
    wire [BITS-1:0] memory_3_scale_8_real_tb;
    wire [BITS-1:0] memory_4_scale_8_real_tb;
    wire [BITS-1:0] memory_5_scale_8_real_tb;
    wire [BITS-1:0] memory_6_scale_8_real_tb;
    wire [BITS-1:0] memory_7_scale_8_real_tb;
    wire [BITS-1:0] memory_8_scale_8_real_tb;
    wire [BITS-1:0] memory_9_scale_8_real_tb;
    wire [BITS-1:0] memory_10_scale_8_real_tb;
    wire [BITS-1:0] memory_11_scale_8_real_tb;
    wire [BITS-1:0] memory_12_scale_8_real_tb;
    wire [BITS-1:0] memory_13_scale_8_real_tb;
    wire [BITS-1:0] memory_14_scale_8_real_tb;
    wire [BITS-1:0] memory_15_scale_8_real_tb;
    wire [BITS-1:0] memory_16_scale_8_real_tb;
    wire [BITS-1:0] memory_17_scale_8_real_tb;
    wire [BITS-1:0] memory_18_scale_8_real_tb;
    wire [BITS-1:0] memory_19_scale_8_real_tb;
    wire [BITS-1:0] memory_20_scale_8_real_tb;
    wire [BITS-1:0] memory_21_scale_8_real_tb;
    wire [BITS-1:0] memory_22_scale_8_real_tb;
    wire [BITS-1:0] memory_23_scale_8_real_tb;
    wire [BITS-1:0] memory_24_scale_8_real_tb;
    wire [BITS-1:0] memory_25_scale_8_real_tb;
    wire [BITS-1:0] memory_26_scale_8_real_tb;
    wire [BITS-1:0] memory_27_scale_8_real_tb;
    wire [BITS-1:0] memory_28_scale_8_real_tb;
    wire [BITS-1:0] memory_29_scale_8_real_tb;
    wire [BITS-1:0] memory_30_scale_8_real_tb;
    wire [BITS-1:0] memory_31_scale_8_real_tb;
    wire [BITS-1:0] memory_0_scale_9_real_tb;
    wire [BITS-1:0] memory_1_scale_9_real_tb;
    wire [BITS-1:0] memory_2_scale_9_real_tb;
    wire [BITS-1:0] memory_3_scale_9_real_tb;
    wire [BITS-1:0] memory_4_scale_9_real_tb;
    wire [BITS-1:0] memory_5_scale_9_real_tb;
    wire [BITS-1:0] memory_6_scale_9_real_tb;
    wire [BITS-1:0] memory_7_scale_9_real_tb;
    wire [BITS-1:0] memory_8_scale_9_real_tb;
    wire [BITS-1:0] memory_9_scale_9_real_tb;
    wire [BITS-1:0] memory_10_scale_9_real_tb;
    wire [BITS-1:0] memory_11_scale_9_real_tb;
    wire [BITS-1:0] memory_12_scale_9_real_tb;
    wire [BITS-1:0] memory_13_scale_9_real_tb;
    wire [BITS-1:0] memory_14_scale_9_real_tb;
    wire [BITS-1:0] memory_15_scale_9_real_tb;
    wire [BITS-1:0] memory_16_scale_9_real_tb;
    wire [BITS-1:0] memory_17_scale_9_real_tb;
    wire [BITS-1:0] memory_18_scale_9_real_tb;
    wire [BITS-1:0] memory_19_scale_9_real_tb;
    wire [BITS-1:0] memory_20_scale_9_real_tb;
    wire [BITS-1:0] memory_21_scale_9_real_tb;
    wire [BITS-1:0] memory_22_scale_9_real_tb;
    wire [BITS-1:0] memory_23_scale_9_real_tb;
    wire [BITS-1:0] memory_24_scale_9_real_tb;
    wire [BITS-1:0] memory_25_scale_9_real_tb;
    wire [BITS-1:0] memory_26_scale_9_real_tb;
    wire [BITS-1:0] memory_27_scale_9_real_tb;
    wire [BITS-1:0] memory_28_scale_9_real_tb;
    wire [BITS-1:0] memory_29_scale_9_real_tb;
    wire [BITS-1:0] memory_30_scale_9_real_tb;
    wire [BITS-1:0] memory_31_scale_9_real_tb;
    wire [BITS-1:0] memory_0_scale_10_real_tb;
    wire [BITS-1:0] memory_1_scale_10_real_tb;
    wire [BITS-1:0] memory_2_scale_10_real_tb;
    wire [BITS-1:0] memory_3_scale_10_real_tb;
    wire [BITS-1:0] memory_4_scale_10_real_tb;
    wire [BITS-1:0] memory_5_scale_10_real_tb;
    wire [BITS-1:0] memory_6_scale_10_real_tb;
    wire [BITS-1:0] memory_7_scale_10_real_tb;
    wire [BITS-1:0] memory_8_scale_10_real_tb;
    wire [BITS-1:0] memory_9_scale_10_real_tb;
    wire [BITS-1:0] memory_10_scale_10_real_tb;
    wire [BITS-1:0] memory_11_scale_10_real_tb;
    wire [BITS-1:0] memory_12_scale_10_real_tb;
    wire [BITS-1:0] memory_13_scale_10_real_tb;
    wire [BITS-1:0] memory_14_scale_10_real_tb;
    wire [BITS-1:0] memory_15_scale_10_real_tb;
    wire [BITS-1:0] memory_16_scale_10_real_tb;
    wire [BITS-1:0] memory_17_scale_10_real_tb;
    wire [BITS-1:0] memory_18_scale_10_real_tb;
    wire [BITS-1:0] memory_19_scale_10_real_tb;
    wire [BITS-1:0] memory_20_scale_10_real_tb;
    wire [BITS-1:0] memory_21_scale_10_real_tb;
    wire [BITS-1:0] memory_22_scale_10_real_tb;
    wire [BITS-1:0] memory_23_scale_10_real_tb;
    wire [BITS-1:0] memory_24_scale_10_real_tb;
    wire [BITS-1:0] memory_25_scale_10_real_tb;
    wire [BITS-1:0] memory_26_scale_10_real_tb;
    wire [BITS-1:0] memory_27_scale_10_real_tb;
    wire [BITS-1:0] memory_28_scale_10_real_tb;
    wire [BITS-1:0] memory_29_scale_10_real_tb;
    wire [BITS-1:0] memory_30_scale_10_real_tb;
    wire [BITS-1:0] memory_31_scale_10_real_tb;
    wire [BITS-1:0] memory_0_scale_11_real_tb;
    wire [BITS-1:0] memory_1_scale_11_real_tb;
    wire [BITS-1:0] memory_2_scale_11_real_tb;
    wire [BITS-1:0] memory_3_scale_11_real_tb;
    wire [BITS-1:0] memory_4_scale_11_real_tb;
    wire [BITS-1:0] memory_5_scale_11_real_tb;
    wire [BITS-1:0] memory_6_scale_11_real_tb;
    wire [BITS-1:0] memory_7_scale_11_real_tb;
    wire [BITS-1:0] memory_8_scale_11_real_tb;
    wire [BITS-1:0] memory_9_scale_11_real_tb;
    wire [BITS-1:0] memory_10_scale_11_real_tb;
    wire [BITS-1:0] memory_11_scale_11_real_tb;
    wire [BITS-1:0] memory_12_scale_11_real_tb;
    wire [BITS-1:0] memory_13_scale_11_real_tb;
    wire [BITS-1:0] memory_14_scale_11_real_tb;
    wire [BITS-1:0] memory_15_scale_11_real_tb;
    wire [BITS-1:0] memory_16_scale_11_real_tb;
    wire [BITS-1:0] memory_17_scale_11_real_tb;
    wire [BITS-1:0] memory_18_scale_11_real_tb;
    wire [BITS-1:0] memory_19_scale_11_real_tb;
    wire [BITS-1:0] memory_20_scale_11_real_tb;
    wire [BITS-1:0] memory_21_scale_11_real_tb;
    wire [BITS-1:0] memory_22_scale_11_real_tb;
    wire [BITS-1:0] memory_23_scale_11_real_tb;
    wire [BITS-1:0] memory_24_scale_11_real_tb;
    wire [BITS-1:0] memory_25_scale_11_real_tb;
    wire [BITS-1:0] memory_26_scale_11_real_tb;
    wire [BITS-1:0] memory_27_scale_11_real_tb;
    wire [BITS-1:0] memory_28_scale_11_real_tb;
    wire [BITS-1:0] memory_29_scale_11_real_tb;
    wire [BITS-1:0] memory_30_scale_11_real_tb;
    wire [BITS-1:0] memory_31_scale_11_real_tb;
    wire [BITS-1:0] memory_0_scale_12_real_tb;
    wire [BITS-1:0] memory_1_scale_12_real_tb;
    wire [BITS-1:0] memory_2_scale_12_real_tb;
    wire [BITS-1:0] memory_3_scale_12_real_tb;
    wire [BITS-1:0] memory_4_scale_12_real_tb;
    wire [BITS-1:0] memory_5_scale_12_real_tb;
    wire [BITS-1:0] memory_6_scale_12_real_tb;
    wire [BITS-1:0] memory_7_scale_12_real_tb;
    wire [BITS-1:0] memory_8_scale_12_real_tb;
    wire [BITS-1:0] memory_9_scale_12_real_tb;
    wire [BITS-1:0] memory_10_scale_12_real_tb;
    wire [BITS-1:0] memory_11_scale_12_real_tb;
    wire [BITS-1:0] memory_12_scale_12_real_tb;
    wire [BITS-1:0] memory_13_scale_12_real_tb;
    wire [BITS-1:0] memory_14_scale_12_real_tb;
    wire [BITS-1:0] memory_15_scale_12_real_tb;
    wire [BITS-1:0] memory_16_scale_12_real_tb;
    wire [BITS-1:0] memory_17_scale_12_real_tb;
    wire [BITS-1:0] memory_18_scale_12_real_tb;
    wire [BITS-1:0] memory_19_scale_12_real_tb;
    wire [BITS-1:0] memory_20_scale_12_real_tb;
    wire [BITS-1:0] memory_21_scale_12_real_tb;
    wire [BITS-1:0] memory_22_scale_12_real_tb;
    wire [BITS-1:0] memory_23_scale_12_real_tb;
    wire [BITS-1:0] memory_24_scale_12_real_tb;
    wire [BITS-1:0] memory_25_scale_12_real_tb;
    wire [BITS-1:0] memory_26_scale_12_real_tb;
    wire [BITS-1:0] memory_27_scale_12_real_tb;
    wire [BITS-1:0] memory_28_scale_12_real_tb;
    wire [BITS-1:0] memory_29_scale_12_real_tb;
    wire [BITS-1:0] memory_30_scale_12_real_tb;
    wire [BITS-1:0] memory_31_scale_12_real_tb;
    wire [BITS-1:0] memory_0_scale_13_real_tb;
    wire [BITS-1:0] memory_1_scale_13_real_tb;
    wire [BITS-1:0] memory_2_scale_13_real_tb;
    wire [BITS-1:0] memory_3_scale_13_real_tb;
    wire [BITS-1:0] memory_4_scale_13_real_tb;
    wire [BITS-1:0] memory_5_scale_13_real_tb;
    wire [BITS-1:0] memory_6_scale_13_real_tb;
    wire [BITS-1:0] memory_7_scale_13_real_tb;
    wire [BITS-1:0] memory_8_scale_13_real_tb;
    wire [BITS-1:0] memory_9_scale_13_real_tb;
    wire [BITS-1:0] memory_10_scale_13_real_tb;
    wire [BITS-1:0] memory_11_scale_13_real_tb;
    wire [BITS-1:0] memory_12_scale_13_real_tb;
    wire [BITS-1:0] memory_13_scale_13_real_tb;
    wire [BITS-1:0] memory_14_scale_13_real_tb;
    wire [BITS-1:0] memory_15_scale_13_real_tb;
    wire [BITS-1:0] memory_16_scale_13_real_tb;
    wire [BITS-1:0] memory_17_scale_13_real_tb;
    wire [BITS-1:0] memory_18_scale_13_real_tb;
    wire [BITS-1:0] memory_19_scale_13_real_tb;
    wire [BITS-1:0] memory_20_scale_13_real_tb;
    wire [BITS-1:0] memory_21_scale_13_real_tb;
    wire [BITS-1:0] memory_22_scale_13_real_tb;
    wire [BITS-1:0] memory_23_scale_13_real_tb;
    wire [BITS-1:0] memory_24_scale_13_real_tb;
    wire [BITS-1:0] memory_25_scale_13_real_tb;
    wire [BITS-1:0] memory_26_scale_13_real_tb;
    wire [BITS-1:0] memory_27_scale_13_real_tb;
    wire [BITS-1:0] memory_28_scale_13_real_tb;
    wire [BITS-1:0] memory_29_scale_13_real_tb;
    wire [BITS-1:0] memory_30_scale_13_real_tb;
    wire [BITS-1:0] memory_31_scale_13_real_tb;
    wire [BITS-1:0] memory_0_scale_14_real_tb;
    wire [BITS-1:0] memory_1_scale_14_real_tb;
    wire [BITS-1:0] memory_2_scale_14_real_tb;
    wire [BITS-1:0] memory_3_scale_14_real_tb;
    wire [BITS-1:0] memory_4_scale_14_real_tb;
    wire [BITS-1:0] memory_5_scale_14_real_tb;
    wire [BITS-1:0] memory_6_scale_14_real_tb;
    wire [BITS-1:0] memory_7_scale_14_real_tb;
    wire [BITS-1:0] memory_8_scale_14_real_tb;
    wire [BITS-1:0] memory_9_scale_14_real_tb;
    wire [BITS-1:0] memory_10_scale_14_real_tb;
    wire [BITS-1:0] memory_11_scale_14_real_tb;
    wire [BITS-1:0] memory_12_scale_14_real_tb;
    wire [BITS-1:0] memory_13_scale_14_real_tb;
    wire [BITS-1:0] memory_14_scale_14_real_tb;
    wire [BITS-1:0] memory_15_scale_14_real_tb;
    wire [BITS-1:0] memory_16_scale_14_real_tb;
    wire [BITS-1:0] memory_17_scale_14_real_tb;
    wire [BITS-1:0] memory_18_scale_14_real_tb;
    wire [BITS-1:0] memory_19_scale_14_real_tb;
    wire [BITS-1:0] memory_20_scale_14_real_tb;
    wire [BITS-1:0] memory_21_scale_14_real_tb;
    wire [BITS-1:0] memory_22_scale_14_real_tb;
    wire [BITS-1:0] memory_23_scale_14_real_tb;
    wire [BITS-1:0] memory_24_scale_14_real_tb;
    wire [BITS-1:0] memory_25_scale_14_real_tb;
    wire [BITS-1:0] memory_26_scale_14_real_tb;
    wire [BITS-1:0] memory_27_scale_14_real_tb;
    wire [BITS-1:0] memory_28_scale_14_real_tb;
    wire [BITS-1:0] memory_29_scale_14_real_tb;
    wire [BITS-1:0] memory_30_scale_14_real_tb;
    wire [BITS-1:0] memory_31_scale_14_real_tb;
    wire [BITS-1:0] memory_0_scale_15_real_tb;
    wire [BITS-1:0] memory_1_scale_15_real_tb;
    wire [BITS-1:0] memory_2_scale_15_real_tb;
    wire [BITS-1:0] memory_3_scale_15_real_tb;
    wire [BITS-1:0] memory_4_scale_15_real_tb;
    wire [BITS-1:0] memory_5_scale_15_real_tb;
    wire [BITS-1:0] memory_6_scale_15_real_tb;
    wire [BITS-1:0] memory_7_scale_15_real_tb;
    wire [BITS-1:0] memory_8_scale_15_real_tb;
    wire [BITS-1:0] memory_9_scale_15_real_tb;
    wire [BITS-1:0] memory_10_scale_15_real_tb;
    wire [BITS-1:0] memory_11_scale_15_real_tb;
    wire [BITS-1:0] memory_12_scale_15_real_tb;
    wire [BITS-1:0] memory_13_scale_15_real_tb;
    wire [BITS-1:0] memory_14_scale_15_real_tb;
    wire [BITS-1:0] memory_15_scale_15_real_tb;
    wire [BITS-1:0] memory_16_scale_15_real_tb;
    wire [BITS-1:0] memory_17_scale_15_real_tb;
    wire [BITS-1:0] memory_18_scale_15_real_tb;
    wire [BITS-1:0] memory_19_scale_15_real_tb;
    wire [BITS-1:0] memory_20_scale_15_real_tb;
    wire [BITS-1:0] memory_21_scale_15_real_tb;
    wire [BITS-1:0] memory_22_scale_15_real_tb;
    wire [BITS-1:0] memory_23_scale_15_real_tb;
    wire [BITS-1:0] memory_24_scale_15_real_tb;
    wire [BITS-1:0] memory_25_scale_15_real_tb;
    wire [BITS-1:0] memory_26_scale_15_real_tb;
    wire [BITS-1:0] memory_27_scale_15_real_tb;
    wire [BITS-1:0] memory_28_scale_15_real_tb;
    wire [BITS-1:0] memory_29_scale_15_real_tb;
    wire [BITS-1:0] memory_30_scale_15_real_tb;
    wire [BITS-1:0] memory_31_scale_15_real_tb;




    wire [BITS-1:0] memory_0_scale_1_imag_tb ;
    wire [BITS-1:0] memory_1_scale_1_imag_tb ;
    wire [BITS-1:0] memory_2_scale_1_imag_tb ;
    wire [BITS-1:0] memory_3_scale_1_imag_tb ;
    wire [BITS-1:0] memory_4_scale_1_imag_tb ;
    wire [BITS-1:0] memory_5_scale_1_imag_tb ;
    wire [BITS-1:0] memory_6_scale_1_imag_tb ;
    wire [BITS-1:0] memory_7_scale_1_imag_tb ;
    wire [BITS-1:0] memory_8_scale_1_imag_tb ;
    wire [BITS-1:0] memory_9_scale_1_imag_tb ;
    wire [BITS-1:0] memory_10_scale_1_imag_tb ;
    wire [BITS-1:0] memory_11_scale_1_imag_tb ;
    wire [BITS-1:0] memory_12_scale_1_imag_tb ;
    wire [BITS-1:0] memory_13_scale_1_imag_tb ;
    wire [BITS-1:0] memory_14_scale_1_imag_tb ;
    wire [BITS-1:0] memory_15_scale_1_imag_tb ;
    wire [BITS-1:0] memory_16_scale_1_imag_tb ;
    wire [BITS-1:0] memory_17_scale_1_imag_tb ;
    wire [BITS-1:0] memory_18_scale_1_imag_tb ;
    wire [BITS-1:0] memory_19_scale_1_imag_tb ;
    wire [BITS-1:0] memory_20_scale_1_imag_tb ;
    wire [BITS-1:0] memory_21_scale_1_imag_tb ;
    wire [BITS-1:0] memory_22_scale_1_imag_tb ;
    wire [BITS-1:0] memory_23_scale_1_imag_tb ;
    wire [BITS-1:0] memory_24_scale_1_imag_tb ;
    wire [BITS-1:0] memory_25_scale_1_imag_tb ;
    wire [BITS-1:0] memory_26_scale_1_imag_tb ;
    wire [BITS-1:0] memory_27_scale_1_imag_tb ;
    wire [BITS-1:0] memory_28_scale_1_imag_tb ;
    wire [BITS-1:0] memory_29_scale_1_imag_tb ;
    wire [BITS-1:0] memory_30_scale_1_imag_tb ;
    wire [BITS-1:0] memory_31_scale_1_imag_tb ;
    wire [BITS-1:0] memory_0_scale_2_imag_tb ;
    wire [BITS-1:0] memory_1_scale_2_imag_tb ;
    wire [BITS-1:0] memory_2_scale_2_imag_tb ;
    wire [BITS-1:0] memory_3_scale_2_imag_tb ;
    wire [BITS-1:0] memory_4_scale_2_imag_tb ;
    wire [BITS-1:0] memory_5_scale_2_imag_tb ;
    wire [BITS-1:0] memory_6_scale_2_imag_tb ;
    wire [BITS-1:0] memory_7_scale_2_imag_tb ;
    wire [BITS-1:0] memory_8_scale_2_imag_tb ;
    wire [BITS-1:0] memory_9_scale_2_imag_tb ;
    wire [BITS-1:0] memory_10_scale_2_imag_tb ;
    wire [BITS-1:0] memory_11_scale_2_imag_tb ;
    wire [BITS-1:0] memory_12_scale_2_imag_tb ;
    wire [BITS-1:0] memory_13_scale_2_imag_tb ;
    wire [BITS-1:0] memory_14_scale_2_imag_tb ;
    wire [BITS-1:0] memory_15_scale_2_imag_tb ;
    wire [BITS-1:0] memory_16_scale_2_imag_tb ;
    wire [BITS-1:0] memory_17_scale_2_imag_tb ;
    wire [BITS-1:0] memory_18_scale_2_imag_tb ;
    wire [BITS-1:0] memory_19_scale_2_imag_tb ;
    wire [BITS-1:0] memory_20_scale_2_imag_tb ;
    wire [BITS-1:0] memory_21_scale_2_imag_tb ;
    wire [BITS-1:0] memory_22_scale_2_imag_tb ;
    wire [BITS-1:0] memory_23_scale_2_imag_tb ;
    wire [BITS-1:0] memory_24_scale_2_imag_tb ;
    wire [BITS-1:0] memory_25_scale_2_imag_tb ;
    wire [BITS-1:0] memory_26_scale_2_imag_tb ;
    wire [BITS-1:0] memory_27_scale_2_imag_tb ;
    wire [BITS-1:0] memory_28_scale_2_imag_tb ;
    wire [BITS-1:0] memory_29_scale_2_imag_tb ;
    wire [BITS-1:0] memory_30_scale_2_imag_tb ;
    wire [BITS-1:0] memory_31_scale_2_imag_tb ;
    wire [BITS-1:0] memory_0_scale_3_imag_tb ;
    wire [BITS-1:0] memory_1_scale_3_imag_tb ;
    wire [BITS-1:0] memory_2_scale_3_imag_tb ;
    wire [BITS-1:0] memory_3_scale_3_imag_tb ;
    wire [BITS-1:0] memory_4_scale_3_imag_tb ;
    wire [BITS-1:0] memory_5_scale_3_imag_tb ;
    wire [BITS-1:0] memory_6_scale_3_imag_tb ;
    wire [BITS-1:0] memory_7_scale_3_imag_tb ;
    wire [BITS-1:0] memory_8_scale_3_imag_tb ;
    wire [BITS-1:0] memory_9_scale_3_imag_tb ;
    wire [BITS-1:0] memory_10_scale_3_imag_tb ;
    wire [BITS-1:0] memory_11_scale_3_imag_tb ;
    wire [BITS-1:0] memory_12_scale_3_imag_tb ;
    wire [BITS-1:0] memory_13_scale_3_imag_tb ;
    wire [BITS-1:0] memory_14_scale_3_imag_tb ;
    wire [BITS-1:0] memory_15_scale_3_imag_tb ;
    wire [BITS-1:0] memory_16_scale_3_imag_tb ;
    wire [BITS-1:0] memory_17_scale_3_imag_tb ;
    wire [BITS-1:0] memory_18_scale_3_imag_tb ;
    wire [BITS-1:0] memory_19_scale_3_imag_tb ;
    wire [BITS-1:0] memory_20_scale_3_imag_tb ;
    wire [BITS-1:0] memory_21_scale_3_imag_tb ;
    wire [BITS-1:0] memory_22_scale_3_imag_tb ;
    wire [BITS-1:0] memory_23_scale_3_imag_tb ;
    wire [BITS-1:0] memory_24_scale_3_imag_tb ;
    wire [BITS-1:0] memory_25_scale_3_imag_tb ;
    wire [BITS-1:0] memory_26_scale_3_imag_tb ;
    wire [BITS-1:0] memory_27_scale_3_imag_tb ;
    wire [BITS-1:0] memory_28_scale_3_imag_tb ;
    wire [BITS-1:0] memory_29_scale_3_imag_tb ;
    wire [BITS-1:0] memory_30_scale_3_imag_tb ;
    wire [BITS-1:0] memory_31_scale_3_imag_tb ;
    wire [BITS-1:0] memory_0_scale_4_imag_tb ;
    wire [BITS-1:0] memory_1_scale_4_imag_tb ;
    wire [BITS-1:0] memory_2_scale_4_imag_tb ;
    wire [BITS-1:0] memory_3_scale_4_imag_tb ;
    wire [BITS-1:0] memory_4_scale_4_imag_tb ;
    wire [BITS-1:0] memory_5_scale_4_imag_tb ;
    wire [BITS-1:0] memory_6_scale_4_imag_tb ;
    wire [BITS-1:0] memory_7_scale_4_imag_tb ;
    wire [BITS-1:0] memory_8_scale_4_imag_tb ;
    wire [BITS-1:0] memory_9_scale_4_imag_tb ;
    wire [BITS-1:0] memory_10_scale_4_imag_tb ;
    wire [BITS-1:0] memory_11_scale_4_imag_tb ;
    wire [BITS-1:0] memory_12_scale_4_imag_tb ;
    wire [BITS-1:0] memory_13_scale_4_imag_tb ;
    wire [BITS-1:0] memory_14_scale_4_imag_tb ;
    wire [BITS-1:0] memory_15_scale_4_imag_tb ;
    wire [BITS-1:0] memory_16_scale_4_imag_tb ;
    wire [BITS-1:0] memory_17_scale_4_imag_tb ;
    wire [BITS-1:0] memory_18_scale_4_imag_tb ;
    wire [BITS-1:0] memory_19_scale_4_imag_tb ;
    wire [BITS-1:0] memory_20_scale_4_imag_tb ;
    wire [BITS-1:0] memory_21_scale_4_imag_tb ;
    wire [BITS-1:0] memory_22_scale_4_imag_tb ;
    wire [BITS-1:0] memory_23_scale_4_imag_tb ;
    wire [BITS-1:0] memory_24_scale_4_imag_tb ;
    wire [BITS-1:0] memory_25_scale_4_imag_tb ;
    wire [BITS-1:0] memory_26_scale_4_imag_tb ;
    wire [BITS-1:0] memory_27_scale_4_imag_tb ;
    wire [BITS-1:0] memory_28_scale_4_imag_tb ;
    wire [BITS-1:0] memory_29_scale_4_imag_tb ;
    wire [BITS-1:0] memory_30_scale_4_imag_tb ;
    wire [BITS-1:0] memory_31_scale_4_imag_tb ;
    wire [BITS-1:0] memory_0_scale_5_imag_tb ;
    wire [BITS-1:0] memory_1_scale_5_imag_tb ;
    wire [BITS-1:0] memory_2_scale_5_imag_tb ;
    wire [BITS-1:0] memory_3_scale_5_imag_tb ;
    wire [BITS-1:0] memory_4_scale_5_imag_tb ;
    wire [BITS-1:0] memory_5_scale_5_imag_tb ;
    wire [BITS-1:0] memory_6_scale_5_imag_tb ;
    wire [BITS-1:0] memory_7_scale_5_imag_tb ;
    wire [BITS-1:0] memory_8_scale_5_imag_tb ;
    wire [BITS-1:0] memory_9_scale_5_imag_tb ;
    wire [BITS-1:0] memory_10_scale_5_imag_tb ;
    wire [BITS-1:0] memory_11_scale_5_imag_tb ;
    wire [BITS-1:0] memory_12_scale_5_imag_tb ;
    wire [BITS-1:0] memory_13_scale_5_imag_tb ;
    wire [BITS-1:0] memory_14_scale_5_imag_tb ;
    wire [BITS-1:0] memory_15_scale_5_imag_tb ;
    wire [BITS-1:0] memory_16_scale_5_imag_tb ;
    wire [BITS-1:0] memory_17_scale_5_imag_tb ;
    wire [BITS-1:0] memory_18_scale_5_imag_tb ;
    wire [BITS-1:0] memory_19_scale_5_imag_tb ;
    wire [BITS-1:0] memory_20_scale_5_imag_tb ;
    wire [BITS-1:0] memory_21_scale_5_imag_tb ;
    wire [BITS-1:0] memory_22_scale_5_imag_tb ;
    wire [BITS-1:0] memory_23_scale_5_imag_tb ;
    wire [BITS-1:0] memory_24_scale_5_imag_tb ;
    wire [BITS-1:0] memory_25_scale_5_imag_tb ;
    wire [BITS-1:0] memory_26_scale_5_imag_tb ;
    wire [BITS-1:0] memory_27_scale_5_imag_tb ;
    wire [BITS-1:0] memory_28_scale_5_imag_tb ;
    wire [BITS-1:0] memory_29_scale_5_imag_tb ;
    wire [BITS-1:0] memory_30_scale_5_imag_tb ;
    wire [BITS-1:0] memory_31_scale_5_imag_tb ;
    wire [BITS-1:0] memory_0_scale_6_imag_tb ;
    wire [BITS-1:0] memory_1_scale_6_imag_tb ;
    wire [BITS-1:0] memory_2_scale_6_imag_tb ;
    wire [BITS-1:0] memory_3_scale_6_imag_tb ;
    wire [BITS-1:0] memory_4_scale_6_imag_tb ;
    wire [BITS-1:0] memory_5_scale_6_imag_tb ;
    wire [BITS-1:0] memory_6_scale_6_imag_tb ;
    wire [BITS-1:0] memory_7_scale_6_imag_tb ;
    wire [BITS-1:0] memory_8_scale_6_imag_tb ;
    wire [BITS-1:0] memory_9_scale_6_imag_tb ;
    wire [BITS-1:0] memory_10_scale_6_imag_tb ;
    wire [BITS-1:0] memory_11_scale_6_imag_tb ;
    wire [BITS-1:0] memory_12_scale_6_imag_tb ;
    wire [BITS-1:0] memory_13_scale_6_imag_tb ;
    wire [BITS-1:0] memory_14_scale_6_imag_tb ;
    wire [BITS-1:0] memory_15_scale_6_imag_tb ;
    wire [BITS-1:0] memory_16_scale_6_imag_tb ;
    wire [BITS-1:0] memory_17_scale_6_imag_tb ;
    wire [BITS-1:0] memory_18_scale_6_imag_tb ;
    wire [BITS-1:0] memory_19_scale_6_imag_tb ;
    wire [BITS-1:0] memory_20_scale_6_imag_tb ;
    wire [BITS-1:0] memory_21_scale_6_imag_tb ;
    wire [BITS-1:0] memory_22_scale_6_imag_tb ;
    wire [BITS-1:0] memory_23_scale_6_imag_tb ;
    wire [BITS-1:0] memory_24_scale_6_imag_tb ;
    wire [BITS-1:0] memory_25_scale_6_imag_tb ;
    wire [BITS-1:0] memory_26_scale_6_imag_tb ;
    wire [BITS-1:0] memory_27_scale_6_imag_tb ;
    wire [BITS-1:0] memory_28_scale_6_imag_tb ;
    wire [BITS-1:0] memory_29_scale_6_imag_tb ;
    wire [BITS-1:0] memory_30_scale_6_imag_tb ;
    wire [BITS-1:0] memory_31_scale_6_imag_tb ;
    wire [BITS-1:0] memory_0_scale_7_imag_tb ;
    wire [BITS-1:0] memory_1_scale_7_imag_tb ;
    wire [BITS-1:0] memory_2_scale_7_imag_tb ;
    wire [BITS-1:0] memory_3_scale_7_imag_tb ;
    wire [BITS-1:0] memory_4_scale_7_imag_tb ;
    wire [BITS-1:0] memory_5_scale_7_imag_tb ;
    wire [BITS-1:0] memory_6_scale_7_imag_tb ;
    wire [BITS-1:0] memory_7_scale_7_imag_tb ;
    wire [BITS-1:0] memory_8_scale_7_imag_tb ;
    wire [BITS-1:0] memory_9_scale_7_imag_tb ;
    wire [BITS-1:0] memory_10_scale_7_imag_tb ;
    wire [BITS-1:0] memory_11_scale_7_imag_tb ;
    wire [BITS-1:0] memory_12_scale_7_imag_tb ;
    wire [BITS-1:0] memory_13_scale_7_imag_tb ;
    wire [BITS-1:0] memory_14_scale_7_imag_tb ;
    wire [BITS-1:0] memory_15_scale_7_imag_tb ;
    wire [BITS-1:0] memory_16_scale_7_imag_tb ;
    wire [BITS-1:0] memory_17_scale_7_imag_tb ;
    wire [BITS-1:0] memory_18_scale_7_imag_tb ;
    wire [BITS-1:0] memory_19_scale_7_imag_tb ;
    wire [BITS-1:0] memory_20_scale_7_imag_tb ;
    wire [BITS-1:0] memory_21_scale_7_imag_tb ;
    wire [BITS-1:0] memory_22_scale_7_imag_tb ;
    wire [BITS-1:0] memory_23_scale_7_imag_tb ;
    wire [BITS-1:0] memory_24_scale_7_imag_tb ;
    wire [BITS-1:0] memory_25_scale_7_imag_tb ;
    wire [BITS-1:0] memory_26_scale_7_imag_tb ;
    wire [BITS-1:0] memory_27_scale_7_imag_tb ;
    wire [BITS-1:0] memory_28_scale_7_imag_tb ;
    wire [BITS-1:0] memory_29_scale_7_imag_tb ;
    wire [BITS-1:0] memory_30_scale_7_imag_tb ;
    wire [BITS-1:0] memory_31_scale_7_imag_tb ;
    wire [BITS-1:0] memory_0_scale_8_imag_tb ;
    wire [BITS-1:0] memory_1_scale_8_imag_tb ;
    wire [BITS-1:0] memory_2_scale_8_imag_tb ;
    wire [BITS-1:0] memory_3_scale_8_imag_tb ;
    wire [BITS-1:0] memory_4_scale_8_imag_tb ;
    wire [BITS-1:0] memory_5_scale_8_imag_tb ;
    wire [BITS-1:0] memory_6_scale_8_imag_tb ;
    wire [BITS-1:0] memory_7_scale_8_imag_tb ;
    wire [BITS-1:0] memory_8_scale_8_imag_tb ;
    wire [BITS-1:0] memory_9_scale_8_imag_tb ;
    wire [BITS-1:0] memory_10_scale_8_imag_tb ;
    wire [BITS-1:0] memory_11_scale_8_imag_tb ;
    wire [BITS-1:0] memory_12_scale_8_imag_tb ;
    wire [BITS-1:0] memory_13_scale_8_imag_tb ;
    wire [BITS-1:0] memory_14_scale_8_imag_tb ;
    wire [BITS-1:0] memory_15_scale_8_imag_tb ;
    wire [BITS-1:0] memory_16_scale_8_imag_tb ;
    wire [BITS-1:0] memory_17_scale_8_imag_tb ;
    wire [BITS-1:0] memory_18_scale_8_imag_tb ;
    wire [BITS-1:0] memory_19_scale_8_imag_tb ;
    wire [BITS-1:0] memory_20_scale_8_imag_tb ;
    wire [BITS-1:0] memory_21_scale_8_imag_tb ;
    wire [BITS-1:0] memory_22_scale_8_imag_tb ;
    wire [BITS-1:0] memory_23_scale_8_imag_tb ;
    wire [BITS-1:0] memory_24_scale_8_imag_tb ;
    wire [BITS-1:0] memory_25_scale_8_imag_tb ;
    wire [BITS-1:0] memory_26_scale_8_imag_tb ;
    wire [BITS-1:0] memory_27_scale_8_imag_tb ;
    wire [BITS-1:0] memory_28_scale_8_imag_tb ;
    wire [BITS-1:0] memory_29_scale_8_imag_tb ;
    wire [BITS-1:0] memory_30_scale_8_imag_tb ;
    wire [BITS-1:0] memory_31_scale_8_imag_tb ;
    wire [BITS-1:0] memory_0_scale_9_imag_tb ;
    wire [BITS-1:0] memory_1_scale_9_imag_tb ;
    wire [BITS-1:0] memory_2_scale_9_imag_tb ;
    wire [BITS-1:0] memory_3_scale_9_imag_tb ;
    wire [BITS-1:0] memory_4_scale_9_imag_tb ;
    wire [BITS-1:0] memory_5_scale_9_imag_tb ;
    wire [BITS-1:0] memory_6_scale_9_imag_tb ;
    wire [BITS-1:0] memory_7_scale_9_imag_tb ;
    wire [BITS-1:0] memory_8_scale_9_imag_tb ;
    wire [BITS-1:0] memory_9_scale_9_imag_tb ;
    wire [BITS-1:0] memory_10_scale_9_imag_tb ;
    wire [BITS-1:0] memory_11_scale_9_imag_tb ;
    wire [BITS-1:0] memory_12_scale_9_imag_tb ;
    wire [BITS-1:0] memory_13_scale_9_imag_tb ;
    wire [BITS-1:0] memory_14_scale_9_imag_tb ;
    wire [BITS-1:0] memory_15_scale_9_imag_tb ;
    wire [BITS-1:0] memory_16_scale_9_imag_tb ;
    wire [BITS-1:0] memory_17_scale_9_imag_tb ;
    wire [BITS-1:0] memory_18_scale_9_imag_tb ;
    wire [BITS-1:0] memory_19_scale_9_imag_tb ;
    wire [BITS-1:0] memory_20_scale_9_imag_tb ;
    wire [BITS-1:0] memory_21_scale_9_imag_tb ;
    wire [BITS-1:0] memory_22_scale_9_imag_tb ;
    wire [BITS-1:0] memory_23_scale_9_imag_tb ;
    wire [BITS-1:0] memory_24_scale_9_imag_tb ;
    wire [BITS-1:0] memory_25_scale_9_imag_tb ;
    wire [BITS-1:0] memory_26_scale_9_imag_tb ;
    wire [BITS-1:0] memory_27_scale_9_imag_tb ;
    wire [BITS-1:0] memory_28_scale_9_imag_tb ;
    wire [BITS-1:0] memory_29_scale_9_imag_tb ;
    wire [BITS-1:0] memory_30_scale_9_imag_tb ;
    wire [BITS-1:0] memory_31_scale_9_imag_tb ;
    wire [BITS-1:0] memory_0_scale_10_imag_tb ;
    wire [BITS-1:0] memory_1_scale_10_imag_tb ;
    wire [BITS-1:0] memory_2_scale_10_imag_tb ;
    wire [BITS-1:0] memory_3_scale_10_imag_tb ;
    wire [BITS-1:0] memory_4_scale_10_imag_tb ;
    wire [BITS-1:0] memory_5_scale_10_imag_tb ;
    wire [BITS-1:0] memory_6_scale_10_imag_tb ;
    wire [BITS-1:0] memory_7_scale_10_imag_tb ;
    wire [BITS-1:0] memory_8_scale_10_imag_tb ;
    wire [BITS-1:0] memory_9_scale_10_imag_tb ;
    wire [BITS-1:0] memory_10_scale_10_imag_tb ;
    wire [BITS-1:0] memory_11_scale_10_imag_tb ;
    wire [BITS-1:0] memory_12_scale_10_imag_tb ;
    wire [BITS-1:0] memory_13_scale_10_imag_tb ;
    wire [BITS-1:0] memory_14_scale_10_imag_tb ;
    wire [BITS-1:0] memory_15_scale_10_imag_tb ;
    wire [BITS-1:0] memory_16_scale_10_imag_tb ;
    wire [BITS-1:0] memory_17_scale_10_imag_tb ;
    wire [BITS-1:0] memory_18_scale_10_imag_tb ;
    wire [BITS-1:0] memory_19_scale_10_imag_tb ;
    wire [BITS-1:0] memory_20_scale_10_imag_tb ;
    wire [BITS-1:0] memory_21_scale_10_imag_tb ;
    wire [BITS-1:0] memory_22_scale_10_imag_tb ;
    wire [BITS-1:0] memory_23_scale_10_imag_tb ;
    wire [BITS-1:0] memory_24_scale_10_imag_tb ;
    wire [BITS-1:0] memory_25_scale_10_imag_tb ;
    wire [BITS-1:0] memory_26_scale_10_imag_tb ;
    wire [BITS-1:0] memory_27_scale_10_imag_tb ;
    wire [BITS-1:0] memory_28_scale_10_imag_tb ;
    wire [BITS-1:0] memory_29_scale_10_imag_tb ;
    wire [BITS-1:0] memory_30_scale_10_imag_tb ;
    wire [BITS-1:0] memory_31_scale_10_imag_tb ;
    wire [BITS-1:0] memory_0_scale_11_imag_tb ;
    wire [BITS-1:0] memory_1_scale_11_imag_tb ;
    wire [BITS-1:0] memory_2_scale_11_imag_tb ;
    wire [BITS-1:0] memory_3_scale_11_imag_tb ;
    wire [BITS-1:0] memory_4_scale_11_imag_tb ;
    wire [BITS-1:0] memory_5_scale_11_imag_tb ;
    wire [BITS-1:0] memory_6_scale_11_imag_tb ;
    wire [BITS-1:0] memory_7_scale_11_imag_tb ;
    wire [BITS-1:0] memory_8_scale_11_imag_tb ;
    wire [BITS-1:0] memory_9_scale_11_imag_tb ;
    wire [BITS-1:0] memory_10_scale_11_imag_tb ;
    wire [BITS-1:0] memory_11_scale_11_imag_tb ;
    wire [BITS-1:0] memory_12_scale_11_imag_tb ;
    wire [BITS-1:0] memory_13_scale_11_imag_tb ;
    wire [BITS-1:0] memory_14_scale_11_imag_tb ;
    wire [BITS-1:0] memory_15_scale_11_imag_tb ;
    wire [BITS-1:0] memory_16_scale_11_imag_tb ;
    wire [BITS-1:0] memory_17_scale_11_imag_tb ;
    wire [BITS-1:0] memory_18_scale_11_imag_tb ;
    wire [BITS-1:0] memory_19_scale_11_imag_tb ;
    wire [BITS-1:0] memory_20_scale_11_imag_tb ;
    wire [BITS-1:0] memory_21_scale_11_imag_tb ;
    wire [BITS-1:0] memory_22_scale_11_imag_tb ;
    wire [BITS-1:0] memory_23_scale_11_imag_tb ;
    wire [BITS-1:0] memory_24_scale_11_imag_tb ;
    wire [BITS-1:0] memory_25_scale_11_imag_tb ;
    wire [BITS-1:0] memory_26_scale_11_imag_tb ;
    wire [BITS-1:0] memory_27_scale_11_imag_tb ;
    wire [BITS-1:0] memory_28_scale_11_imag_tb ;
    wire [BITS-1:0] memory_29_scale_11_imag_tb ;
    wire [BITS-1:0] memory_30_scale_11_imag_tb ;
    wire [BITS-1:0] memory_31_scale_11_imag_tb ;
    wire [BITS-1:0] memory_0_scale_12_imag_tb ;
    wire [BITS-1:0] memory_1_scale_12_imag_tb ;
    wire [BITS-1:0] memory_2_scale_12_imag_tb ;
    wire [BITS-1:0] memory_3_scale_12_imag_tb ;
    wire [BITS-1:0] memory_4_scale_12_imag_tb ;
    wire [BITS-1:0] memory_5_scale_12_imag_tb ;
    wire [BITS-1:0] memory_6_scale_12_imag_tb ;
    wire [BITS-1:0] memory_7_scale_12_imag_tb ;
    wire [BITS-1:0] memory_8_scale_12_imag_tb ;
    wire [BITS-1:0] memory_9_scale_12_imag_tb ;
    wire [BITS-1:0] memory_10_scale_12_imag_tb ;
    wire [BITS-1:0] memory_11_scale_12_imag_tb ;
    wire [BITS-1:0] memory_12_scale_12_imag_tb ;
    wire [BITS-1:0] memory_13_scale_12_imag_tb ;
    wire [BITS-1:0] memory_14_scale_12_imag_tb ;
    wire [BITS-1:0] memory_15_scale_12_imag_tb ;
    wire [BITS-1:0] memory_16_scale_12_imag_tb ;
    wire [BITS-1:0] memory_17_scale_12_imag_tb ;
    wire [BITS-1:0] memory_18_scale_12_imag_tb ;
    wire [BITS-1:0] memory_19_scale_12_imag_tb ;
    wire [BITS-1:0] memory_20_scale_12_imag_tb ;
    wire [BITS-1:0] memory_21_scale_12_imag_tb ;
    wire [BITS-1:0] memory_22_scale_12_imag_tb ;
    wire [BITS-1:0] memory_23_scale_12_imag_tb ;
    wire [BITS-1:0] memory_24_scale_12_imag_tb ;
    wire [BITS-1:0] memory_25_scale_12_imag_tb ;
    wire [BITS-1:0] memory_26_scale_12_imag_tb ;
    wire [BITS-1:0] memory_27_scale_12_imag_tb ;
    wire [BITS-1:0] memory_28_scale_12_imag_tb ;
    wire [BITS-1:0] memory_29_scale_12_imag_tb ;
    wire [BITS-1:0] memory_30_scale_12_imag_tb ;
    wire [BITS-1:0] memory_31_scale_12_imag_tb ;
    wire [BITS-1:0] memory_0_scale_13_imag_tb ;
    wire [BITS-1:0] memory_1_scale_13_imag_tb ;
    wire [BITS-1:0] memory_2_scale_13_imag_tb ;
    wire [BITS-1:0] memory_3_scale_13_imag_tb ;
    wire [BITS-1:0] memory_4_scale_13_imag_tb ;
    wire [BITS-1:0] memory_5_scale_13_imag_tb ;
    wire [BITS-1:0] memory_6_scale_13_imag_tb ;
    wire [BITS-1:0] memory_7_scale_13_imag_tb ;
    wire [BITS-1:0] memory_8_scale_13_imag_tb ;
    wire [BITS-1:0] memory_9_scale_13_imag_tb ;
    wire [BITS-1:0] memory_10_scale_13_imag_tb ;
    wire [BITS-1:0] memory_11_scale_13_imag_tb ;
    wire [BITS-1:0] memory_12_scale_13_imag_tb ;
    wire [BITS-1:0] memory_13_scale_13_imag_tb ;
    wire [BITS-1:0] memory_14_scale_13_imag_tb ;
    wire [BITS-1:0] memory_15_scale_13_imag_tb ;
    wire [BITS-1:0] memory_16_scale_13_imag_tb ;
    wire [BITS-1:0] memory_17_scale_13_imag_tb ;
    wire [BITS-1:0] memory_18_scale_13_imag_tb ;
    wire [BITS-1:0] memory_19_scale_13_imag_tb ;
    wire [BITS-1:0] memory_20_scale_13_imag_tb ;
    wire [BITS-1:0] memory_21_scale_13_imag_tb ;
    wire [BITS-1:0] memory_22_scale_13_imag_tb ;
    wire [BITS-1:0] memory_23_scale_13_imag_tb ;
    wire [BITS-1:0] memory_24_scale_13_imag_tb ;
    wire [BITS-1:0] memory_25_scale_13_imag_tb ;
    wire [BITS-1:0] memory_26_scale_13_imag_tb ;
    wire [BITS-1:0] memory_27_scale_13_imag_tb ;
    wire [BITS-1:0] memory_28_scale_13_imag_tb ;
    wire [BITS-1:0] memory_29_scale_13_imag_tb ;
    wire [BITS-1:0] memory_30_scale_13_imag_tb ;
    wire [BITS-1:0] memory_31_scale_13_imag_tb ;
    wire [BITS-1:0] memory_0_scale_14_imag_tb ;
    wire [BITS-1:0] memory_1_scale_14_imag_tb ;
    wire [BITS-1:0] memory_2_scale_14_imag_tb ;
    wire [BITS-1:0] memory_3_scale_14_imag_tb ;
    wire [BITS-1:0] memory_4_scale_14_imag_tb ;
    wire [BITS-1:0] memory_5_scale_14_imag_tb ;
    wire [BITS-1:0] memory_6_scale_14_imag_tb ;
    wire [BITS-1:0] memory_7_scale_14_imag_tb ;
    wire [BITS-1:0] memory_8_scale_14_imag_tb ;
    wire [BITS-1:0] memory_9_scale_14_imag_tb ;
    wire [BITS-1:0] memory_10_scale_14_imag_tb ;
    wire [BITS-1:0] memory_11_scale_14_imag_tb ;
    wire [BITS-1:0] memory_12_scale_14_imag_tb ;
    wire [BITS-1:0] memory_13_scale_14_imag_tb ;
    wire [BITS-1:0] memory_14_scale_14_imag_tb ;
    wire [BITS-1:0] memory_15_scale_14_imag_tb ;
    wire [BITS-1:0] memory_16_scale_14_imag_tb ;
    wire [BITS-1:0] memory_17_scale_14_imag_tb ;
    wire [BITS-1:0] memory_18_scale_14_imag_tb ;
    wire [BITS-1:0] memory_19_scale_14_imag_tb ;
    wire [BITS-1:0] memory_20_scale_14_imag_tb ;
    wire [BITS-1:0] memory_21_scale_14_imag_tb ;
    wire [BITS-1:0] memory_22_scale_14_imag_tb ;
    wire [BITS-1:0] memory_23_scale_14_imag_tb ;
    wire [BITS-1:0] memory_24_scale_14_imag_tb ;
    wire [BITS-1:0] memory_25_scale_14_imag_tb ;
    wire [BITS-1:0] memory_26_scale_14_imag_tb ;
    wire [BITS-1:0] memory_27_scale_14_imag_tb ;
    wire [BITS-1:0] memory_28_scale_14_imag_tb ;
    wire [BITS-1:0] memory_29_scale_14_imag_tb ;
    wire [BITS-1:0] memory_30_scale_14_imag_tb ;
    wire [BITS-1:0] memory_31_scale_14_imag_tb ;
    wire [BITS-1:0] memory_0_scale_15_imag_tb ;
    wire [BITS-1:0] memory_1_scale_15_imag_tb ;
    wire [BITS-1:0] memory_2_scale_15_imag_tb ;
    wire [BITS-1:0] memory_3_scale_15_imag_tb ;
    wire [BITS-1:0] memory_4_scale_15_imag_tb ;
    wire [BITS-1:0] memory_5_scale_15_imag_tb ;
    wire [BITS-1:0] memory_6_scale_15_imag_tb ;
    wire [BITS-1:0] memory_7_scale_15_imag_tb ;
    wire [BITS-1:0] memory_8_scale_15_imag_tb ;
    wire [BITS-1:0] memory_9_scale_15_imag_tb ;
    wire [BITS-1:0] memory_10_scale_15_imag_tb ;
    wire [BITS-1:0] memory_11_scale_15_imag_tb ;
    wire [BITS-1:0] memory_12_scale_15_imag_tb ;
    wire [BITS-1:0] memory_13_scale_15_imag_tb ;
    wire [BITS-1:0] memory_14_scale_15_imag_tb ;
    wire [BITS-1:0] memory_15_scale_15_imag_tb ;
    wire [BITS-1:0] memory_16_scale_15_imag_tb ;
    wire [BITS-1:0] memory_17_scale_15_imag_tb ;
    wire [BITS-1:0] memory_18_scale_15_imag_tb ;
    wire [BITS-1:0] memory_19_scale_15_imag_tb ;
    wire [BITS-1:0] memory_20_scale_15_imag_tb ;
    wire [BITS-1:0] memory_21_scale_15_imag_tb ;
    wire [BITS-1:0] memory_22_scale_15_imag_tb ;
    wire [BITS-1:0] memory_23_scale_15_imag_tb ;
    wire [BITS-1:0] memory_24_scale_15_imag_tb ;
    wire [BITS-1:0] memory_25_scale_15_imag_tb ;
    wire [BITS-1:0] memory_26_scale_15_imag_tb ;
    wire [BITS-1:0] memory_27_scale_15_imag_tb ;
    wire [BITS-1:0] memory_28_scale_15_imag_tb ;
    wire [BITS-1:0] memory_29_scale_15_imag_tb ;
    wire [BITS-1:0] memory_30_scale_15_imag_tb ;
    wire [BITS-1:0] memory_31_scale_15_imag_tb ;



    
    cwt_top_module #(.BITS(BITS)) UUT_CWT_TOP
    (
.ready_inputs(ready_inputs_tb) ,
.clk(clk_tb),
.rst(rst_tb),
.read_scale_ram_addresses(read_scale_ram_addresses),
.x0_r(x0_r_tb) ,
.x1_r(x1_r_tb) ,
.x2_r(x2_r_tb) ,
.x3_r(x3_r_tb) ,
.x4_r(x4_r_tb) ,
.x5_r(x5_r_tb) ,
.x6_r(x6_r_tb) ,
.x7_r(x7_r_tb) ,
.x8_r(x8_r_tb) ,
.x9_r(x9_r_tb) ,
.x10_r(x10_r_tb) ,
.x11_r(x11_r_tb) ,
.x12_r(x12_r_tb) ,
.x13_r(x13_r_tb) ,
.x14_r(x14_r_tb) ,
.x15_r(x15_r_tb) ,
.x16_r(x16_r_tb) ,
.x17_r(x17_r_tb) ,
.x18_r(x18_r_tb) ,
.x19_r(x19_r_tb) ,
.x20_r(x20_r_tb) ,
.x21_r(x21_r_tb) ,
.x22_r(x22_r_tb) ,
.x23_r(x23_r_tb) ,
.x24_r(x24_r_tb) ,
.x25_r(x25_r_tb) ,
.x26_r(x26_r_tb) ,
.x27_r(x27_r_tb) ,
.x28_r(x28_r_tb) ,
.x29_r(x29_r_tb) ,
.x30_r(x30_r_tb) ,
.x31_r(x31_r_tb) ,
.x32_r(x32_r_tb) ,
.x33_r(x33_r_tb) ,
.x34_r(x34_r_tb) ,
.x35_r(x35_r_tb) ,
.x36_r(x36_r_tb) ,
.x37_r(x37_r_tb) ,
.x38_r(x38_r_tb) ,
.x39_r(x39_r_tb) ,
.x40_r(x40_r_tb) ,
.x41_r(x41_r_tb) ,
.x42_r(x42_r_tb) ,
.x43_r(x43_r_tb) ,
.x44_r(x44_r_tb) ,
.x45_r(x45_r_tb) ,
.x46_r(x46_r_tb) ,
.x47_r(x47_r_tb) ,
.x48_r(x48_r_tb) ,
.x49_r(x49_r_tb) ,
.x50_r(x50_r_tb) ,
.x51_r(x51_r_tb) ,
.x52_r(x52_r_tb) ,
.x53_r(x53_r_tb) ,
.x54_r(x54_r_tb) ,
.x55_r(x55_r_tb) ,
.x56_r(x56_r_tb) ,
.x57_r(x57_r_tb) ,
.x58_r(x58_r_tb) ,
.x59_r(x59_r_tb) ,
.x60_r(x60_r_tb) ,
.x61_r(x61_r_tb) ,
.x62_r(x62_r_tb) ,
.x63_r(x63_r_tb) ,
.x64_r(x64_r_tb) ,
.x65_r(x65_r_tb) ,
.x66_r(x66_r_tb) ,
.x67_r(x67_r_tb) ,
.x68_r(x68_r_tb) ,
.x69_r(x69_r_tb) ,
.x70_r(x70_r_tb) ,
.x71_r(x71_r_tb) ,
.x72_r(x72_r_tb) ,
.x73_r(x73_r_tb) ,
.x74_r(x74_r_tb) ,
.x75_r(x75_r_tb) ,
.x76_r(x76_r_tb) ,
.x77_r(x77_r_tb) ,
.x78_r(x78_r_tb) ,
.x79_r(x79_r_tb) ,
.x80_r(x80_r_tb) ,
.x81_r(x81_r_tb) ,
.x82_r(x82_r_tb) ,
.x83_r(x83_r_tb) ,
.x84_r(x84_r_tb) ,
.x85_r(x85_r_tb) ,
.x86_r(x86_r_tb) ,
.x87_r(x87_r_tb) ,
.x88_r(x88_r_tb) ,
.x89_r(x89_r_tb) ,
.x90_r(x90_r_tb) ,
.x91_r(x91_r_tb) ,
.x92_r(x92_r_tb) ,
.x93_r(x93_r_tb) ,
.x94_r(x94_r_tb) ,
.x95_r(x95_r_tb) ,
.x96_r(x96_r_tb) ,
.x97_r(x97_r_tb) ,
.x98_r(x98_r_tb) ,
.x99_r(x99_r_tb) ,
.x100_r(x100_r_tb) ,
.x101_r(x101_r_tb) ,
.x102_r(x102_r_tb) ,
.x103_r(x103_r_tb) ,
.x104_r(x104_r_tb) ,
.x105_r(x105_r_tb) ,
.x106_r(x106_r_tb) ,
.x107_r(x107_r_tb) ,
.x108_r(x108_r_tb) ,
.x109_r(x109_r_tb) ,
.x110_r(x110_r_tb) ,
.x111_r(x111_r_tb) ,
.x112_r(x112_r_tb) ,
.x113_r(x113_r_tb) ,
.x114_r(x114_r_tb) ,
.x115_r(x115_r_tb) ,
.x116_r(x116_r_tb) ,
.x117_r(x117_r_tb) ,
.x118_r(x118_r_tb) ,
.x119_r(x119_r_tb) ,
.x120_r(x120_r_tb) ,
.x121_r(x121_r_tb) ,
.x122_r(x122_r_tb) ,
.x123_r(x123_r_tb) ,
.x124_r(x124_r_tb) ,
.x125_r(x125_r_tb) ,
.x126_r(x126_r_tb) ,
.x127_r(x127_r_tb) ,
.memory_0_scale_1_real(memory_0_scale_1_real_tb),
.memory_1_scale_1_real(memory_1_scale_1_real_tb),
.memory_2_scale_1_real(memory_2_scale_1_real_tb),
.memory_3_scale_1_real(memory_3_scale_1_real_tb),
.memory_4_scale_1_real(memory_4_scale_1_real_tb),
.memory_5_scale_1_real(memory_5_scale_1_real_tb),
.memory_6_scale_1_real(memory_6_scale_1_real_tb),
.memory_7_scale_1_real(memory_7_scale_1_real_tb),
.memory_8_scale_1_real(memory_8_scale_1_real_tb),
.memory_9_scale_1_real(memory_9_scale_1_real_tb),
.memory_10_scale_1_real(memory_10_scale_1_real_tb),
.memory_11_scale_1_real(memory_11_scale_1_real_tb),
.memory_12_scale_1_real(memory_12_scale_1_real_tb),
.memory_13_scale_1_real(memory_13_scale_1_real_tb),
.memory_14_scale_1_real(memory_14_scale_1_real_tb),
.memory_15_scale_1_real(memory_15_scale_1_real_tb),
.memory_16_scale_1_real(memory_16_scale_1_real_tb),
.memory_17_scale_1_real(memory_17_scale_1_real_tb),
.memory_18_scale_1_real(memory_18_scale_1_real_tb),
.memory_19_scale_1_real(memory_19_scale_1_real_tb),
.memory_20_scale_1_real(memory_20_scale_1_real_tb),
.memory_21_scale_1_real(memory_21_scale_1_real_tb),
.memory_22_scale_1_real(memory_22_scale_1_real_tb),
.memory_23_scale_1_real(memory_23_scale_1_real_tb),
.memory_24_scale_1_real(memory_24_scale_1_real_tb),
.memory_25_scale_1_real(memory_25_scale_1_real_tb),
.memory_26_scale_1_real(memory_26_scale_1_real_tb),
.memory_27_scale_1_real(memory_27_scale_1_real_tb),
.memory_28_scale_1_real(memory_28_scale_1_real_tb),
.memory_29_scale_1_real(memory_29_scale_1_real_tb),
.memory_30_scale_1_real(memory_30_scale_1_real_tb),
.memory_31_scale_1_real(memory_31_scale_1_real_tb),
.memory_0_scale_2_real(memory_0_scale_2_real_tb),
.memory_1_scale_2_real(memory_1_scale_2_real_tb),
.memory_2_scale_2_real(memory_2_scale_2_real_tb),
.memory_3_scale_2_real(memory_3_scale_2_real_tb),
.memory_4_scale_2_real(memory_4_scale_2_real_tb),
.memory_5_scale_2_real(memory_5_scale_2_real_tb),
.memory_6_scale_2_real(memory_6_scale_2_real_tb),
.memory_7_scale_2_real(memory_7_scale_2_real_tb),
.memory_8_scale_2_real(memory_8_scale_2_real_tb),
.memory_9_scale_2_real(memory_9_scale_2_real_tb),
.memory_10_scale_2_real(memory_10_scale_2_real_tb),
.memory_11_scale_2_real(memory_11_scale_2_real_tb),
.memory_12_scale_2_real(memory_12_scale_2_real_tb),
.memory_13_scale_2_real(memory_13_scale_2_real_tb),
.memory_14_scale_2_real(memory_14_scale_2_real_tb),
.memory_15_scale_2_real(memory_15_scale_2_real_tb),
.memory_16_scale_2_real(memory_16_scale_2_real_tb),
.memory_17_scale_2_real(memory_17_scale_2_real_tb),
.memory_18_scale_2_real(memory_18_scale_2_real_tb),
.memory_19_scale_2_real(memory_19_scale_2_real_tb),
.memory_20_scale_2_real(memory_20_scale_2_real_tb),
.memory_21_scale_2_real(memory_21_scale_2_real_tb),
.memory_22_scale_2_real(memory_22_scale_2_real_tb),
.memory_23_scale_2_real(memory_23_scale_2_real_tb),
.memory_24_scale_2_real(memory_24_scale_2_real_tb),
.memory_25_scale_2_real(memory_25_scale_2_real_tb),
.memory_26_scale_2_real(memory_26_scale_2_real_tb),
.memory_27_scale_2_real(memory_27_scale_2_real_tb),
.memory_28_scale_2_real(memory_28_scale_2_real_tb),
.memory_29_scale_2_real(memory_29_scale_2_real_tb),
.memory_30_scale_2_real(memory_30_scale_2_real_tb),
.memory_31_scale_2_real(memory_31_scale_2_real_tb),
.memory_0_scale_3_real(memory_0_scale_3_real_tb),
.memory_1_scale_3_real(memory_1_scale_3_real_tb),
.memory_2_scale_3_real(memory_2_scale_3_real_tb),
.memory_3_scale_3_real(memory_3_scale_3_real_tb),
.memory_4_scale_3_real(memory_4_scale_3_real_tb),
.memory_5_scale_3_real(memory_5_scale_3_real_tb),
.memory_6_scale_3_real(memory_6_scale_3_real_tb),
.memory_7_scale_3_real(memory_7_scale_3_real_tb),
.memory_8_scale_3_real(memory_8_scale_3_real_tb),
.memory_9_scale_3_real(memory_9_scale_3_real_tb),
.memory_10_scale_3_real(memory_10_scale_3_real_tb),
.memory_11_scale_3_real(memory_11_scale_3_real_tb),
.memory_12_scale_3_real(memory_12_scale_3_real_tb),
.memory_13_scale_3_real(memory_13_scale_3_real_tb),
.memory_14_scale_3_real(memory_14_scale_3_real_tb),
.memory_15_scale_3_real(memory_15_scale_3_real_tb),
.memory_16_scale_3_real(memory_16_scale_3_real_tb),
.memory_17_scale_3_real(memory_17_scale_3_real_tb),
.memory_18_scale_3_real(memory_18_scale_3_real_tb),
.memory_19_scale_3_real(memory_19_scale_3_real_tb),
.memory_20_scale_3_real(memory_20_scale_3_real_tb),
.memory_21_scale_3_real(memory_21_scale_3_real_tb),
.memory_22_scale_3_real(memory_22_scale_3_real_tb),
.memory_23_scale_3_real(memory_23_scale_3_real_tb),
.memory_24_scale_3_real(memory_24_scale_3_real_tb),
.memory_25_scale_3_real(memory_25_scale_3_real_tb),
.memory_26_scale_3_real(memory_26_scale_3_real_tb),
.memory_27_scale_3_real(memory_27_scale_3_real_tb),
.memory_28_scale_3_real(memory_28_scale_3_real_tb),
.memory_29_scale_3_real(memory_29_scale_3_real_tb),
.memory_30_scale_3_real(memory_30_scale_3_real_tb),
.memory_31_scale_3_real(memory_31_scale_3_real_tb),
.memory_0_scale_4_real(memory_0_scale_4_real_tb),
.memory_1_scale_4_real(memory_1_scale_4_real_tb),
.memory_2_scale_4_real(memory_2_scale_4_real_tb),
.memory_3_scale_4_real(memory_3_scale_4_real_tb),
.memory_4_scale_4_real(memory_4_scale_4_real_tb),
.memory_5_scale_4_real(memory_5_scale_4_real_tb),
.memory_6_scale_4_real(memory_6_scale_4_real_tb),
.memory_7_scale_4_real(memory_7_scale_4_real_tb),
.memory_8_scale_4_real(memory_8_scale_4_real_tb),
.memory_9_scale_4_real(memory_9_scale_4_real_tb),
.memory_10_scale_4_real(memory_10_scale_4_real_tb),
.memory_11_scale_4_real(memory_11_scale_4_real_tb),
.memory_12_scale_4_real(memory_12_scale_4_real_tb),
.memory_13_scale_4_real(memory_13_scale_4_real_tb),
.memory_14_scale_4_real(memory_14_scale_4_real_tb),
.memory_15_scale_4_real(memory_15_scale_4_real_tb),
.memory_16_scale_4_real(memory_16_scale_4_real_tb),
.memory_17_scale_4_real(memory_17_scale_4_real_tb),
.memory_18_scale_4_real(memory_18_scale_4_real_tb),
.memory_19_scale_4_real(memory_19_scale_4_real_tb),
.memory_20_scale_4_real(memory_20_scale_4_real_tb),
.memory_21_scale_4_real(memory_21_scale_4_real_tb),
.memory_22_scale_4_real(memory_22_scale_4_real_tb),
.memory_23_scale_4_real(memory_23_scale_4_real_tb),
.memory_24_scale_4_real(memory_24_scale_4_real_tb),
.memory_25_scale_4_real(memory_25_scale_4_real_tb),
.memory_26_scale_4_real(memory_26_scale_4_real_tb),
.memory_27_scale_4_real(memory_27_scale_4_real_tb),
.memory_28_scale_4_real(memory_28_scale_4_real_tb),
.memory_29_scale_4_real(memory_29_scale_4_real_tb),
.memory_30_scale_4_real(memory_30_scale_4_real_tb),
.memory_31_scale_4_real(memory_31_scale_4_real_tb),
.memory_0_scale_5_real(memory_0_scale_5_real_tb),
.memory_1_scale_5_real(memory_1_scale_5_real_tb),
.memory_2_scale_5_real(memory_2_scale_5_real_tb),
.memory_3_scale_5_real(memory_3_scale_5_real_tb),
.memory_4_scale_5_real(memory_4_scale_5_real_tb),
.memory_5_scale_5_real(memory_5_scale_5_real_tb),
.memory_6_scale_5_real(memory_6_scale_5_real_tb),
.memory_7_scale_5_real(memory_7_scale_5_real_tb),
.memory_8_scale_5_real(memory_8_scale_5_real_tb),
.memory_9_scale_5_real(memory_9_scale_5_real_tb),
.memory_10_scale_5_real(memory_10_scale_5_real_tb),
.memory_11_scale_5_real(memory_11_scale_5_real_tb),
.memory_12_scale_5_real(memory_12_scale_5_real_tb),
.memory_13_scale_5_real(memory_13_scale_5_real_tb),
.memory_14_scale_5_real(memory_14_scale_5_real_tb),
.memory_15_scale_5_real(memory_15_scale_5_real_tb),
.memory_16_scale_5_real(memory_16_scale_5_real_tb),
.memory_17_scale_5_real(memory_17_scale_5_real_tb),
.memory_18_scale_5_real(memory_18_scale_5_real_tb),
.memory_19_scale_5_real(memory_19_scale_5_real_tb),
.memory_20_scale_5_real(memory_20_scale_5_real_tb),
.memory_21_scale_5_real(memory_21_scale_5_real_tb),
.memory_22_scale_5_real(memory_22_scale_5_real_tb),
.memory_23_scale_5_real(memory_23_scale_5_real_tb),
.memory_24_scale_5_real(memory_24_scale_5_real_tb),
.memory_25_scale_5_real(memory_25_scale_5_real_tb),
.memory_26_scale_5_real(memory_26_scale_5_real_tb),
.memory_27_scale_5_real(memory_27_scale_5_real_tb),
.memory_28_scale_5_real(memory_28_scale_5_real_tb),
.memory_29_scale_5_real(memory_29_scale_5_real_tb),
.memory_30_scale_5_real(memory_30_scale_5_real_tb),
.memory_31_scale_5_real(memory_31_scale_5_real_tb),
.memory_0_scale_6_real(memory_0_scale_6_real_tb),
.memory_1_scale_6_real(memory_1_scale_6_real_tb),
.memory_2_scale_6_real(memory_2_scale_6_real_tb),
.memory_3_scale_6_real(memory_3_scale_6_real_tb),
.memory_4_scale_6_real(memory_4_scale_6_real_tb),
.memory_5_scale_6_real(memory_5_scale_6_real_tb),
.memory_6_scale_6_real(memory_6_scale_6_real_tb),
.memory_7_scale_6_real(memory_7_scale_6_real_tb),
.memory_8_scale_6_real(memory_8_scale_6_real_tb),
.memory_9_scale_6_real(memory_9_scale_6_real_tb),
.memory_10_scale_6_real(memory_10_scale_6_real_tb),
.memory_11_scale_6_real(memory_11_scale_6_real_tb),
.memory_12_scale_6_real(memory_12_scale_6_real_tb),
.memory_13_scale_6_real(memory_13_scale_6_real_tb),
.memory_14_scale_6_real(memory_14_scale_6_real_tb),
.memory_15_scale_6_real(memory_15_scale_6_real_tb),
.memory_16_scale_6_real(memory_16_scale_6_real_tb),
.memory_17_scale_6_real(memory_17_scale_6_real_tb),
.memory_18_scale_6_real(memory_18_scale_6_real_tb),
.memory_19_scale_6_real(memory_19_scale_6_real_tb),
.memory_20_scale_6_real(memory_20_scale_6_real_tb),
.memory_21_scale_6_real(memory_21_scale_6_real_tb),
.memory_22_scale_6_real(memory_22_scale_6_real_tb),
.memory_23_scale_6_real(memory_23_scale_6_real_tb),
.memory_24_scale_6_real(memory_24_scale_6_real_tb),
.memory_25_scale_6_real(memory_25_scale_6_real_tb),
.memory_26_scale_6_real(memory_26_scale_6_real_tb),
.memory_27_scale_6_real(memory_27_scale_6_real_tb),
.memory_28_scale_6_real(memory_28_scale_6_real_tb),
.memory_29_scale_6_real(memory_29_scale_6_real_tb),
.memory_30_scale_6_real(memory_30_scale_6_real_tb),
.memory_31_scale_6_real(memory_31_scale_6_real_tb),
.memory_0_scale_7_real(memory_0_scale_7_real_tb),
.memory_1_scale_7_real(memory_1_scale_7_real_tb),
.memory_2_scale_7_real(memory_2_scale_7_real_tb),
.memory_3_scale_7_real(memory_3_scale_7_real_tb),
.memory_4_scale_7_real(memory_4_scale_7_real_tb),
.memory_5_scale_7_real(memory_5_scale_7_real_tb),
.memory_6_scale_7_real(memory_6_scale_7_real_tb),
.memory_7_scale_7_real(memory_7_scale_7_real_tb),
.memory_8_scale_7_real(memory_8_scale_7_real_tb),
.memory_9_scale_7_real(memory_9_scale_7_real_tb),
.memory_10_scale_7_real(memory_10_scale_7_real_tb),
.memory_11_scale_7_real(memory_11_scale_7_real_tb),
.memory_12_scale_7_real(memory_12_scale_7_real_tb),
.memory_13_scale_7_real(memory_13_scale_7_real_tb),
.memory_14_scale_7_real(memory_14_scale_7_real_tb),
.memory_15_scale_7_real(memory_15_scale_7_real_tb),
.memory_16_scale_7_real(memory_16_scale_7_real_tb),
.memory_17_scale_7_real(memory_17_scale_7_real_tb),
.memory_18_scale_7_real(memory_18_scale_7_real_tb),
.memory_19_scale_7_real(memory_19_scale_7_real_tb),
.memory_20_scale_7_real(memory_20_scale_7_real_tb),
.memory_21_scale_7_real(memory_21_scale_7_real_tb),
.memory_22_scale_7_real(memory_22_scale_7_real_tb),
.memory_23_scale_7_real(memory_23_scale_7_real_tb),
.memory_24_scale_7_real(memory_24_scale_7_real_tb),
.memory_25_scale_7_real(memory_25_scale_7_real_tb),
.memory_26_scale_7_real(memory_26_scale_7_real_tb),
.memory_27_scale_7_real(memory_27_scale_7_real_tb),
.memory_28_scale_7_real(memory_28_scale_7_real_tb),
.memory_29_scale_7_real(memory_29_scale_7_real_tb),
.memory_30_scale_7_real(memory_30_scale_7_real_tb),
.memory_31_scale_7_real(memory_31_scale_7_real_tb),
.memory_0_scale_8_real(memory_0_scale_8_real_tb),
.memory_1_scale_8_real(memory_1_scale_8_real_tb),
.memory_2_scale_8_real(memory_2_scale_8_real_tb),
.memory_3_scale_8_real(memory_3_scale_8_real_tb),
.memory_4_scale_8_real(memory_4_scale_8_real_tb),
.memory_5_scale_8_real(memory_5_scale_8_real_tb),
.memory_6_scale_8_real(memory_6_scale_8_real_tb),
.memory_7_scale_8_real(memory_7_scale_8_real_tb),
.memory_8_scale_8_real(memory_8_scale_8_real_tb),
.memory_9_scale_8_real(memory_9_scale_8_real_tb),
.memory_10_scale_8_real(memory_10_scale_8_real_tb),
.memory_11_scale_8_real(memory_11_scale_8_real_tb),
.memory_12_scale_8_real(memory_12_scale_8_real_tb),
.memory_13_scale_8_real(memory_13_scale_8_real_tb),
.memory_14_scale_8_real(memory_14_scale_8_real_tb),
.memory_15_scale_8_real(memory_15_scale_8_real_tb),
.memory_16_scale_8_real(memory_16_scale_8_real_tb),
.memory_17_scale_8_real(memory_17_scale_8_real_tb),
.memory_18_scale_8_real(memory_18_scale_8_real_tb),
.memory_19_scale_8_real(memory_19_scale_8_real_tb),
.memory_20_scale_8_real(memory_20_scale_8_real_tb),
.memory_21_scale_8_real(memory_21_scale_8_real_tb),
.memory_22_scale_8_real(memory_22_scale_8_real_tb),
.memory_23_scale_8_real(memory_23_scale_8_real_tb),
.memory_24_scale_8_real(memory_24_scale_8_real_tb),
.memory_25_scale_8_real(memory_25_scale_8_real_tb),
.memory_26_scale_8_real(memory_26_scale_8_real_tb),
.memory_27_scale_8_real(memory_27_scale_8_real_tb),
.memory_28_scale_8_real(memory_28_scale_8_real_tb),
.memory_29_scale_8_real(memory_29_scale_8_real_tb),
.memory_30_scale_8_real(memory_30_scale_8_real_tb),
.memory_31_scale_8_real(memory_31_scale_8_real_tb),
.memory_0_scale_9_real(memory_0_scale_9_real_tb),
.memory_1_scale_9_real(memory_1_scale_9_real_tb),
.memory_2_scale_9_real(memory_2_scale_9_real_tb),
.memory_3_scale_9_real(memory_3_scale_9_real_tb),
.memory_4_scale_9_real(memory_4_scale_9_real_tb),
.memory_5_scale_9_real(memory_5_scale_9_real_tb),
.memory_6_scale_9_real(memory_6_scale_9_real_tb),
.memory_7_scale_9_real(memory_7_scale_9_real_tb),
.memory_8_scale_9_real(memory_8_scale_9_real_tb),
.memory_9_scale_9_real(memory_9_scale_9_real_tb),
.memory_10_scale_9_real(memory_10_scale_9_real_tb),
.memory_11_scale_9_real(memory_11_scale_9_real_tb),
.memory_12_scale_9_real(memory_12_scale_9_real_tb),
.memory_13_scale_9_real(memory_13_scale_9_real_tb),
.memory_14_scale_9_real(memory_14_scale_9_real_tb),
.memory_15_scale_9_real(memory_15_scale_9_real_tb),
.memory_16_scale_9_real(memory_16_scale_9_real_tb),
.memory_17_scale_9_real(memory_17_scale_9_real_tb),
.memory_18_scale_9_real(memory_18_scale_9_real_tb),
.memory_19_scale_9_real(memory_19_scale_9_real_tb),
.memory_20_scale_9_real(memory_20_scale_9_real_tb),
.memory_21_scale_9_real(memory_21_scale_9_real_tb),
.memory_22_scale_9_real(memory_22_scale_9_real_tb),
.memory_23_scale_9_real(memory_23_scale_9_real_tb),
.memory_24_scale_9_real(memory_24_scale_9_real_tb),
.memory_25_scale_9_real(memory_25_scale_9_real_tb),
.memory_26_scale_9_real(memory_26_scale_9_real_tb),
.memory_27_scale_9_real(memory_27_scale_9_real_tb),
.memory_28_scale_9_real(memory_28_scale_9_real_tb),
.memory_29_scale_9_real(memory_29_scale_9_real_tb),
.memory_30_scale_9_real(memory_30_scale_9_real_tb),
.memory_31_scale_9_real(memory_31_scale_9_real_tb),
.memory_0_scale_10_real(memory_0_scale_10_real_tb),
.memory_1_scale_10_real(memory_1_scale_10_real_tb),
.memory_2_scale_10_real(memory_2_scale_10_real_tb),
.memory_3_scale_10_real(memory_3_scale_10_real_tb),
.memory_4_scale_10_real(memory_4_scale_10_real_tb),
.memory_5_scale_10_real(memory_5_scale_10_real_tb),
.memory_6_scale_10_real(memory_6_scale_10_real_tb),
.memory_7_scale_10_real(memory_7_scale_10_real_tb),
.memory_8_scale_10_real(memory_8_scale_10_real_tb),
.memory_9_scale_10_real(memory_9_scale_10_real_tb),
.memory_10_scale_10_real(memory_10_scale_10_real_tb),
.memory_11_scale_10_real(memory_11_scale_10_real_tb),
.memory_12_scale_10_real(memory_12_scale_10_real_tb),
.memory_13_scale_10_real(memory_13_scale_10_real_tb),
.memory_14_scale_10_real(memory_14_scale_10_real_tb),
.memory_15_scale_10_real(memory_15_scale_10_real_tb),
.memory_16_scale_10_real(memory_16_scale_10_real_tb),
.memory_17_scale_10_real(memory_17_scale_10_real_tb),
.memory_18_scale_10_real(memory_18_scale_10_real_tb),
.memory_19_scale_10_real(memory_19_scale_10_real_tb),
.memory_20_scale_10_real(memory_20_scale_10_real_tb),
.memory_21_scale_10_real(memory_21_scale_10_real_tb),
.memory_22_scale_10_real(memory_22_scale_10_real_tb),
.memory_23_scale_10_real(memory_23_scale_10_real_tb),
.memory_24_scale_10_real(memory_24_scale_10_real_tb),
.memory_25_scale_10_real(memory_25_scale_10_real_tb),
.memory_26_scale_10_real(memory_26_scale_10_real_tb),
.memory_27_scale_10_real(memory_27_scale_10_real_tb),
.memory_28_scale_10_real(memory_28_scale_10_real_tb),
.memory_29_scale_10_real(memory_29_scale_10_real_tb),
.memory_30_scale_10_real(memory_30_scale_10_real_tb),
.memory_31_scale_10_real(memory_31_scale_10_real_tb),
.memory_0_scale_11_real(memory_0_scale_11_real_tb),
.memory_1_scale_11_real(memory_1_scale_11_real_tb),
.memory_2_scale_11_real(memory_2_scale_11_real_tb),
.memory_3_scale_11_real(memory_3_scale_11_real_tb),
.memory_4_scale_11_real(memory_4_scale_11_real_tb),
.memory_5_scale_11_real(memory_5_scale_11_real_tb),
.memory_6_scale_11_real(memory_6_scale_11_real_tb),
.memory_7_scale_11_real(memory_7_scale_11_real_tb),
.memory_8_scale_11_real(memory_8_scale_11_real_tb),
.memory_9_scale_11_real(memory_9_scale_11_real_tb),
.memory_10_scale_11_real(memory_10_scale_11_real_tb),
.memory_11_scale_11_real(memory_11_scale_11_real_tb),
.memory_12_scale_11_real(memory_12_scale_11_real_tb),
.memory_13_scale_11_real(memory_13_scale_11_real_tb),
.memory_14_scale_11_real(memory_14_scale_11_real_tb),
.memory_15_scale_11_real(memory_15_scale_11_real_tb),
.memory_16_scale_11_real(memory_16_scale_11_real_tb),
.memory_17_scale_11_real(memory_17_scale_11_real_tb),
.memory_18_scale_11_real(memory_18_scale_11_real_tb),
.memory_19_scale_11_real(memory_19_scale_11_real_tb),
.memory_20_scale_11_real(memory_20_scale_11_real_tb),
.memory_21_scale_11_real(memory_21_scale_11_real_tb),
.memory_22_scale_11_real(memory_22_scale_11_real_tb),
.memory_23_scale_11_real(memory_23_scale_11_real_tb),
.memory_24_scale_11_real(memory_24_scale_11_real_tb),
.memory_25_scale_11_real(memory_25_scale_11_real_tb),
.memory_26_scale_11_real(memory_26_scale_11_real_tb),
.memory_27_scale_11_real(memory_27_scale_11_real_tb),
.memory_28_scale_11_real(memory_28_scale_11_real_tb),
.memory_29_scale_11_real(memory_29_scale_11_real_tb),
.memory_30_scale_11_real(memory_30_scale_11_real_tb),
.memory_31_scale_11_real(memory_31_scale_11_real_tb),
.memory_0_scale_12_real(memory_0_scale_12_real_tb),
.memory_1_scale_12_real(memory_1_scale_12_real_tb),
.memory_2_scale_12_real(memory_2_scale_12_real_tb),
.memory_3_scale_12_real(memory_3_scale_12_real_tb),
.memory_4_scale_12_real(memory_4_scale_12_real_tb),
.memory_5_scale_12_real(memory_5_scale_12_real_tb),
.memory_6_scale_12_real(memory_6_scale_12_real_tb),
.memory_7_scale_12_real(memory_7_scale_12_real_tb),
.memory_8_scale_12_real(memory_8_scale_12_real_tb),
.memory_9_scale_12_real(memory_9_scale_12_real_tb),
.memory_10_scale_12_real(memory_10_scale_12_real_tb),
.memory_11_scale_12_real(memory_11_scale_12_real_tb),
.memory_12_scale_12_real(memory_12_scale_12_real_tb),
.memory_13_scale_12_real(memory_13_scale_12_real_tb),
.memory_14_scale_12_real(memory_14_scale_12_real_tb),
.memory_15_scale_12_real(memory_15_scale_12_real_tb),
.memory_16_scale_12_real(memory_16_scale_12_real_tb),
.memory_17_scale_12_real(memory_17_scale_12_real_tb),
.memory_18_scale_12_real(memory_18_scale_12_real_tb),
.memory_19_scale_12_real(memory_19_scale_12_real_tb),
.memory_20_scale_12_real(memory_20_scale_12_real_tb),
.memory_21_scale_12_real(memory_21_scale_12_real_tb),
.memory_22_scale_12_real(memory_22_scale_12_real_tb),
.memory_23_scale_12_real(memory_23_scale_12_real_tb),
.memory_24_scale_12_real(memory_24_scale_12_real_tb),
.memory_25_scale_12_real(memory_25_scale_12_real_tb),
.memory_26_scale_12_real(memory_26_scale_12_real_tb),
.memory_27_scale_12_real(memory_27_scale_12_real_tb),
.memory_28_scale_12_real(memory_28_scale_12_real_tb),
.memory_29_scale_12_real(memory_29_scale_12_real_tb),
.memory_30_scale_12_real(memory_30_scale_12_real_tb),
.memory_31_scale_12_real(memory_31_scale_12_real_tb),
.memory_0_scale_13_real(memory_0_scale_13_real_tb),
.memory_1_scale_13_real(memory_1_scale_13_real_tb),
.memory_2_scale_13_real(memory_2_scale_13_real_tb),
.memory_3_scale_13_real(memory_3_scale_13_real_tb),
.memory_4_scale_13_real(memory_4_scale_13_real_tb),
.memory_5_scale_13_real(memory_5_scale_13_real_tb),
.memory_6_scale_13_real(memory_6_scale_13_real_tb),
.memory_7_scale_13_real(memory_7_scale_13_real_tb),
.memory_8_scale_13_real(memory_8_scale_13_real_tb),
.memory_9_scale_13_real(memory_9_scale_13_real_tb),
.memory_10_scale_13_real(memory_10_scale_13_real_tb),
.memory_11_scale_13_real(memory_11_scale_13_real_tb),
.memory_12_scale_13_real(memory_12_scale_13_real_tb),
.memory_13_scale_13_real(memory_13_scale_13_real_tb),
.memory_14_scale_13_real(memory_14_scale_13_real_tb),
.memory_15_scale_13_real(memory_15_scale_13_real_tb),
.memory_16_scale_13_real(memory_16_scale_13_real_tb),
.memory_17_scale_13_real(memory_17_scale_13_real_tb),
.memory_18_scale_13_real(memory_18_scale_13_real_tb),
.memory_19_scale_13_real(memory_19_scale_13_real_tb),
.memory_20_scale_13_real(memory_20_scale_13_real_tb),
.memory_21_scale_13_real(memory_21_scale_13_real_tb),
.memory_22_scale_13_real(memory_22_scale_13_real_tb),
.memory_23_scale_13_real(memory_23_scale_13_real_tb),
.memory_24_scale_13_real(memory_24_scale_13_real_tb),
.memory_25_scale_13_real(memory_25_scale_13_real_tb),
.memory_26_scale_13_real(memory_26_scale_13_real_tb),
.memory_27_scale_13_real(memory_27_scale_13_real_tb),
.memory_28_scale_13_real(memory_28_scale_13_real_tb),
.memory_29_scale_13_real(memory_29_scale_13_real_tb),
.memory_30_scale_13_real(memory_30_scale_13_real_tb),
.memory_31_scale_13_real(memory_31_scale_13_real_tb),
.memory_0_scale_14_real(memory_0_scale_14_real_tb),
.memory_1_scale_14_real(memory_1_scale_14_real_tb),
.memory_2_scale_14_real(memory_2_scale_14_real_tb),
.memory_3_scale_14_real(memory_3_scale_14_real_tb),
.memory_4_scale_14_real(memory_4_scale_14_real_tb),
.memory_5_scale_14_real(memory_5_scale_14_real_tb),
.memory_6_scale_14_real(memory_6_scale_14_real_tb),
.memory_7_scale_14_real(memory_7_scale_14_real_tb),
.memory_8_scale_14_real(memory_8_scale_14_real_tb),
.memory_9_scale_14_real(memory_9_scale_14_real_tb),
.memory_10_scale_14_real(memory_10_scale_14_real_tb),
.memory_11_scale_14_real(memory_11_scale_14_real_tb),
.memory_12_scale_14_real(memory_12_scale_14_real_tb),
.memory_13_scale_14_real(memory_13_scale_14_real_tb),
.memory_14_scale_14_real(memory_14_scale_14_real_tb),
.memory_15_scale_14_real(memory_15_scale_14_real_tb),
.memory_16_scale_14_real(memory_16_scale_14_real_tb),
.memory_17_scale_14_real(memory_17_scale_14_real_tb),
.memory_18_scale_14_real(memory_18_scale_14_real_tb),
.memory_19_scale_14_real(memory_19_scale_14_real_tb),
.memory_20_scale_14_real(memory_20_scale_14_real_tb),
.memory_21_scale_14_real(memory_21_scale_14_real_tb),
.memory_22_scale_14_real(memory_22_scale_14_real_tb),
.memory_23_scale_14_real(memory_23_scale_14_real_tb),
.memory_24_scale_14_real(memory_24_scale_14_real_tb),
.memory_25_scale_14_real(memory_25_scale_14_real_tb),
.memory_26_scale_14_real(memory_26_scale_14_real_tb),
.memory_27_scale_14_real(memory_27_scale_14_real_tb),
.memory_28_scale_14_real(memory_28_scale_14_real_tb),
.memory_29_scale_14_real(memory_29_scale_14_real_tb),
.memory_30_scale_14_real(memory_30_scale_14_real_tb),
.memory_31_scale_14_real(memory_31_scale_14_real_tb),
.memory_0_scale_15_real(memory_0_scale_15_real_tb),
.memory_1_scale_15_real(memory_1_scale_15_real_tb),
.memory_2_scale_15_real(memory_2_scale_15_real_tb),
.memory_3_scale_15_real(memory_3_scale_15_real_tb),
.memory_4_scale_15_real(memory_4_scale_15_real_tb),
.memory_5_scale_15_real(memory_5_scale_15_real_tb),
.memory_6_scale_15_real(memory_6_scale_15_real_tb),
.memory_7_scale_15_real(memory_7_scale_15_real_tb),
.memory_8_scale_15_real(memory_8_scale_15_real_tb),
.memory_9_scale_15_real(memory_9_scale_15_real_tb),
.memory_10_scale_15_real(memory_10_scale_15_real_tb),
.memory_11_scale_15_real(memory_11_scale_15_real_tb),
.memory_12_scale_15_real(memory_12_scale_15_real_tb),
.memory_13_scale_15_real(memory_13_scale_15_real_tb),
.memory_14_scale_15_real(memory_14_scale_15_real_tb),
.memory_15_scale_15_real(memory_15_scale_15_real_tb),
.memory_16_scale_15_real(memory_16_scale_15_real_tb),
.memory_17_scale_15_real(memory_17_scale_15_real_tb),
.memory_18_scale_15_real(memory_18_scale_15_real_tb),
.memory_19_scale_15_real(memory_19_scale_15_real_tb),
.memory_20_scale_15_real(memory_20_scale_15_real_tb),
.memory_21_scale_15_real(memory_21_scale_15_real_tb),
.memory_22_scale_15_real(memory_22_scale_15_real_tb),
.memory_23_scale_15_real(memory_23_scale_15_real_tb),
.memory_24_scale_15_real(memory_24_scale_15_real_tb),
.memory_25_scale_15_real(memory_25_scale_15_real_tb),
.memory_26_scale_15_real(memory_26_scale_15_real_tb),
.memory_27_scale_15_real(memory_27_scale_15_real_tb),
.memory_28_scale_15_real(memory_28_scale_15_real_tb),
.memory_29_scale_15_real(memory_29_scale_15_real_tb),
.memory_30_scale_15_real(memory_30_scale_15_real_tb),
.memory_31_scale_15_real(memory_31_scale_15_real_tb),





.x0_i(x0_i_tb) ,
.x1_i(x1_i_tb) ,
.x2_i(x2_i_tb) ,
.x3_i(x3_i_tb) ,
.x4_i(x4_i_tb) ,
.x5_i(x5_i_tb) ,
.x6_i(x6_i_tb) ,
.x7_i(x7_i_tb) ,
.x8_i(x8_i_tb) ,
.x9_i(x9_i_tb) ,
.x10_i(x10_i_tb) ,
.x11_i(x11_i_tb) ,
.x12_i(x12_i_tb) ,
.x13_i(x13_i_tb) ,
.x14_i(x14_i_tb) ,
.x15_i(x15_i_tb) ,
.x16_i(x16_i_tb) ,
.x17_i(x17_i_tb) ,
.x18_i(x18_i_tb) ,
.x19_i(x19_i_tb) ,
.x20_i(x20_i_tb) ,
.x21_i(x21_i_tb) ,
.x22_i(x22_i_tb) ,
.x23_i(x23_i_tb) ,
.x24_i(x24_i_tb) ,
.x25_i(x25_i_tb) ,
.x26_i(x26_i_tb) ,
.x27_i(x27_i_tb) ,
.x28_i(x28_i_tb) ,
.x29_i(x29_i_tb) ,
.x30_i(x30_i_tb) ,
.x31_i(x31_i_tb) ,
.x32_i(x32_i_tb) ,
.x33_i(x33_i_tb) ,
.x34_i(x34_i_tb) ,
.x35_i(x35_i_tb) ,
.x36_i(x36_i_tb) ,
.x37_i(x37_i_tb) ,
.x38_i(x38_i_tb) ,
.x39_i(x39_i_tb) ,
.x40_i(x40_i_tb) ,
.x41_i(x41_i_tb) ,
.x42_i(x42_i_tb) ,
.x43_i(x43_i_tb) ,
.x44_i(x44_i_tb) ,
.x45_i(x45_i_tb) ,
.x46_i(x46_i_tb) ,
.x47_i(x47_i_tb) ,
.x48_i(x48_i_tb) ,
.x49_i(x49_i_tb) ,
.x50_i(x50_i_tb) ,
.x51_i(x51_i_tb) ,
.x52_i(x52_i_tb) ,
.x53_i(x53_i_tb) ,
.x54_i(x54_i_tb) ,
.x55_i(x55_i_tb) ,
.x56_i(x56_i_tb) ,
.x57_i(x57_i_tb) ,
.x58_i(x58_i_tb) ,
.x59_i(x59_i_tb) ,
.x60_i(x60_i_tb) ,
.x61_i(x61_i_tb) ,
.x62_i(x62_i_tb) ,
.x63_i(x63_i_tb) ,
.x64_i(x64_i_tb) ,
.x65_i(x65_i_tb) ,
.x66_i(x66_i_tb) ,
.x67_i(x67_i_tb) ,
.x68_i(x68_i_tb) ,
.x69_i(x69_i_tb) ,
.x70_i(x70_i_tb) ,
.x71_i(x71_i_tb) ,
.x72_i(x72_i_tb) ,
.x73_i(x73_i_tb) ,
.x74_i(x74_i_tb) ,
.x75_i(x75_i_tb) ,
.x76_i(x76_i_tb) ,
.x77_i(x77_i_tb) ,
.x78_i(x78_i_tb) ,
.x79_i(x79_i_tb) ,
.x80_i(x80_i_tb) ,
.x81_i(x81_i_tb) ,
.x82_i(x82_i_tb) ,
.x83_i(x83_i_tb) ,
.x84_i(x84_i_tb) ,
.x85_i(x85_i_tb) ,
.x86_i(x86_i_tb) ,
.x87_i(x87_i_tb) ,
.x88_i(x88_i_tb) ,
.x89_i(x89_i_tb) ,
.x90_i(x90_i_tb) ,
.x91_i(x91_i_tb) ,
.x92_i(x92_i_tb) ,
.x93_i(x93_i_tb) ,
.x94_i(x94_i_tb) ,
.x95_i(x95_i_tb) ,
.x96_i(x96_i_tb) ,
.x97_i(x97_i_tb) ,
.x98_i(x98_i_tb) ,
.x99_i(x99_i_tb) ,
.x100_i(x100_i_tb) ,
.x101_i(x101_i_tb) ,
.x102_i(x102_i_tb) ,
.x103_i(x103_i_tb) ,
.x104_i(x104_i_tb) ,
.x105_i(x105_i_tb) ,
.x106_i(x106_i_tb) ,
.x107_i(x107_i_tb) ,
.x108_i(x108_i_tb) ,
.x109_i(x109_i_tb) ,
.x110_i(x110_i_tb) ,
.x111_i(x111_i_tb) ,
.x112_i(x112_i_tb) ,
.x113_i(x113_i_tb) ,
.x114_i(x114_i_tb) ,
.x115_i(x115_i_tb) ,
.x116_i(x116_i_tb) ,
.x117_i(x117_i_tb) ,
.x118_i(x118_i_tb) ,
.x119_i(x119_i_tb) ,
.x120_i(x120_i_tb) ,
.x121_i(x121_i_tb) ,
.x122_i(x122_i_tb) ,
.x123_i(x123_i_tb) ,
.x124_i(x124_i_tb) ,
.x125_i(x125_i_tb) ,
.x126_i(x126_i_tb) ,
.x127_i(x127_i_tb) ,
.memory_0_scale_1_imag(memory_0_scale_1_imag_tb),
.memory_1_scale_1_imag(memory_1_scale_1_imag_tb),
.memory_2_scale_1_imag(memory_2_scale_1_imag_tb),
.memory_3_scale_1_imag(memory_3_scale_1_imag_tb),
.memory_4_scale_1_imag(memory_4_scale_1_imag_tb),
.memory_5_scale_1_imag(memory_5_scale_1_imag_tb),
.memory_6_scale_1_imag(memory_6_scale_1_imag_tb),
.memory_7_scale_1_imag(memory_7_scale_1_imag_tb),
.memory_8_scale_1_imag(memory_8_scale_1_imag_tb),
.memory_9_scale_1_imag(memory_9_scale_1_imag_tb),
.memory_10_scale_1_imag(memory_10_scale_1_imag_tb),
.memory_11_scale_1_imag(memory_11_scale_1_imag_tb),
.memory_12_scale_1_imag(memory_12_scale_1_imag_tb),
.memory_13_scale_1_imag(memory_13_scale_1_imag_tb),
.memory_14_scale_1_imag(memory_14_scale_1_imag_tb),
.memory_15_scale_1_imag(memory_15_scale_1_imag_tb),
.memory_16_scale_1_imag(memory_16_scale_1_imag_tb),
.memory_17_scale_1_imag(memory_17_scale_1_imag_tb),
.memory_18_scale_1_imag(memory_18_scale_1_imag_tb),
.memory_19_scale_1_imag(memory_19_scale_1_imag_tb),
.memory_20_scale_1_imag(memory_20_scale_1_imag_tb),
.memory_21_scale_1_imag(memory_21_scale_1_imag_tb),
.memory_22_scale_1_imag(memory_22_scale_1_imag_tb),
.memory_23_scale_1_imag(memory_23_scale_1_imag_tb),
.memory_24_scale_1_imag(memory_24_scale_1_imag_tb),
.memory_25_scale_1_imag(memory_25_scale_1_imag_tb),
.memory_26_scale_1_imag(memory_26_scale_1_imag_tb),
.memory_27_scale_1_imag(memory_27_scale_1_imag_tb),
.memory_28_scale_1_imag(memory_28_scale_1_imag_tb),
.memory_29_scale_1_imag(memory_29_scale_1_imag_tb),
.memory_30_scale_1_imag(memory_30_scale_1_imag_tb),
.memory_31_scale_1_imag(memory_31_scale_1_imag_tb),
.memory_0_scale_2_imag(memory_0_scale_2_imag_tb),
.memory_1_scale_2_imag(memory_1_scale_2_imag_tb),
.memory_2_scale_2_imag(memory_2_scale_2_imag_tb),
.memory_3_scale_2_imag(memory_3_scale_2_imag_tb),
.memory_4_scale_2_imag(memory_4_scale_2_imag_tb),
.memory_5_scale_2_imag(memory_5_scale_2_imag_tb),
.memory_6_scale_2_imag(memory_6_scale_2_imag_tb),
.memory_7_scale_2_imag(memory_7_scale_2_imag_tb),
.memory_8_scale_2_imag(memory_8_scale_2_imag_tb),
.memory_9_scale_2_imag(memory_9_scale_2_imag_tb),
.memory_10_scale_2_imag(memory_10_scale_2_imag_tb),
.memory_11_scale_2_imag(memory_11_scale_2_imag_tb),
.memory_12_scale_2_imag(memory_12_scale_2_imag_tb),
.memory_13_scale_2_imag(memory_13_scale_2_imag_tb),
.memory_14_scale_2_imag(memory_14_scale_2_imag_tb),
.memory_15_scale_2_imag(memory_15_scale_2_imag_tb),
.memory_16_scale_2_imag(memory_16_scale_2_imag_tb),
.memory_17_scale_2_imag(memory_17_scale_2_imag_tb),
.memory_18_scale_2_imag(memory_18_scale_2_imag_tb),
.memory_19_scale_2_imag(memory_19_scale_2_imag_tb),
.memory_20_scale_2_imag(memory_20_scale_2_imag_tb),
.memory_21_scale_2_imag(memory_21_scale_2_imag_tb),
.memory_22_scale_2_imag(memory_22_scale_2_imag_tb),
.memory_23_scale_2_imag(memory_23_scale_2_imag_tb),
.memory_24_scale_2_imag(memory_24_scale_2_imag_tb),
.memory_25_scale_2_imag(memory_25_scale_2_imag_tb),
.memory_26_scale_2_imag(memory_26_scale_2_imag_tb),
.memory_27_scale_2_imag(memory_27_scale_2_imag_tb),
.memory_28_scale_2_imag(memory_28_scale_2_imag_tb),
.memory_29_scale_2_imag(memory_29_scale_2_imag_tb),
.memory_30_scale_2_imag(memory_30_scale_2_imag_tb),
.memory_31_scale_2_imag(memory_31_scale_2_imag_tb),
.memory_0_scale_3_imag(memory_0_scale_3_imag_tb),
.memory_1_scale_3_imag(memory_1_scale_3_imag_tb),
.memory_2_scale_3_imag(memory_2_scale_3_imag_tb),
.memory_3_scale_3_imag(memory_3_scale_3_imag_tb),
.memory_4_scale_3_imag(memory_4_scale_3_imag_tb),
.memory_5_scale_3_imag(memory_5_scale_3_imag_tb),
.memory_6_scale_3_imag(memory_6_scale_3_imag_tb),
.memory_7_scale_3_imag(memory_7_scale_3_imag_tb),
.memory_8_scale_3_imag(memory_8_scale_3_imag_tb),
.memory_9_scale_3_imag(memory_9_scale_3_imag_tb),
.memory_10_scale_3_imag(memory_10_scale_3_imag_tb),
.memory_11_scale_3_imag(memory_11_scale_3_imag_tb),
.memory_12_scale_3_imag(memory_12_scale_3_imag_tb),
.memory_13_scale_3_imag(memory_13_scale_3_imag_tb),
.memory_14_scale_3_imag(memory_14_scale_3_imag_tb),
.memory_15_scale_3_imag(memory_15_scale_3_imag_tb),
.memory_16_scale_3_imag(memory_16_scale_3_imag_tb),
.memory_17_scale_3_imag(memory_17_scale_3_imag_tb),
.memory_18_scale_3_imag(memory_18_scale_3_imag_tb),
.memory_19_scale_3_imag(memory_19_scale_3_imag_tb),
.memory_20_scale_3_imag(memory_20_scale_3_imag_tb),
.memory_21_scale_3_imag(memory_21_scale_3_imag_tb),
.memory_22_scale_3_imag(memory_22_scale_3_imag_tb),
.memory_23_scale_3_imag(memory_23_scale_3_imag_tb),
.memory_24_scale_3_imag(memory_24_scale_3_imag_tb),
.memory_25_scale_3_imag(memory_25_scale_3_imag_tb),
.memory_26_scale_3_imag(memory_26_scale_3_imag_tb),
.memory_27_scale_3_imag(memory_27_scale_3_imag_tb),
.memory_28_scale_3_imag(memory_28_scale_3_imag_tb),
.memory_29_scale_3_imag(memory_29_scale_3_imag_tb),
.memory_30_scale_3_imag(memory_30_scale_3_imag_tb),
.memory_31_scale_3_imag(memory_31_scale_3_imag_tb),
.memory_0_scale_4_imag(memory_0_scale_4_imag_tb),
.memory_1_scale_4_imag(memory_1_scale_4_imag_tb),
.memory_2_scale_4_imag(memory_2_scale_4_imag_tb),
.memory_3_scale_4_imag(memory_3_scale_4_imag_tb),
.memory_4_scale_4_imag(memory_4_scale_4_imag_tb),
.memory_5_scale_4_imag(memory_5_scale_4_imag_tb),
.memory_6_scale_4_imag(memory_6_scale_4_imag_tb),
.memory_7_scale_4_imag(memory_7_scale_4_imag_tb),
.memory_8_scale_4_imag(memory_8_scale_4_imag_tb),
.memory_9_scale_4_imag(memory_9_scale_4_imag_tb),
.memory_10_scale_4_imag(memory_10_scale_4_imag_tb),
.memory_11_scale_4_imag(memory_11_scale_4_imag_tb),
.memory_12_scale_4_imag(memory_12_scale_4_imag_tb),
.memory_13_scale_4_imag(memory_13_scale_4_imag_tb),
.memory_14_scale_4_imag(memory_14_scale_4_imag_tb),
.memory_15_scale_4_imag(memory_15_scale_4_imag_tb),
.memory_16_scale_4_imag(memory_16_scale_4_imag_tb),
.memory_17_scale_4_imag(memory_17_scale_4_imag_tb),
.memory_18_scale_4_imag(memory_18_scale_4_imag_tb),
.memory_19_scale_4_imag(memory_19_scale_4_imag_tb),
.memory_20_scale_4_imag(memory_20_scale_4_imag_tb),
.memory_21_scale_4_imag(memory_21_scale_4_imag_tb),
.memory_22_scale_4_imag(memory_22_scale_4_imag_tb),
.memory_23_scale_4_imag(memory_23_scale_4_imag_tb),
.memory_24_scale_4_imag(memory_24_scale_4_imag_tb),
.memory_25_scale_4_imag(memory_25_scale_4_imag_tb),
.memory_26_scale_4_imag(memory_26_scale_4_imag_tb),
.memory_27_scale_4_imag(memory_27_scale_4_imag_tb),
.memory_28_scale_4_imag(memory_28_scale_4_imag_tb),
.memory_29_scale_4_imag(memory_29_scale_4_imag_tb),
.memory_30_scale_4_imag(memory_30_scale_4_imag_tb),
.memory_31_scale_4_imag(memory_31_scale_4_imag_tb),
.memory_0_scale_5_imag(memory_0_scale_5_imag_tb),
.memory_1_scale_5_imag(memory_1_scale_5_imag_tb),
.memory_2_scale_5_imag(memory_2_scale_5_imag_tb),
.memory_3_scale_5_imag(memory_3_scale_5_imag_tb),
.memory_4_scale_5_imag(memory_4_scale_5_imag_tb),
.memory_5_scale_5_imag(memory_5_scale_5_imag_tb),
.memory_6_scale_5_imag(memory_6_scale_5_imag_tb),
.memory_7_scale_5_imag(memory_7_scale_5_imag_tb),
.memory_8_scale_5_imag(memory_8_scale_5_imag_tb),
.memory_9_scale_5_imag(memory_9_scale_5_imag_tb),
.memory_10_scale_5_imag(memory_10_scale_5_imag_tb),
.memory_11_scale_5_imag(memory_11_scale_5_imag_tb),
.memory_12_scale_5_imag(memory_12_scale_5_imag_tb),
.memory_13_scale_5_imag(memory_13_scale_5_imag_tb),
.memory_14_scale_5_imag(memory_14_scale_5_imag_tb),
.memory_15_scale_5_imag(memory_15_scale_5_imag_tb),
.memory_16_scale_5_imag(memory_16_scale_5_imag_tb),
.memory_17_scale_5_imag(memory_17_scale_5_imag_tb),
.memory_18_scale_5_imag(memory_18_scale_5_imag_tb),
.memory_19_scale_5_imag(memory_19_scale_5_imag_tb),
.memory_20_scale_5_imag(memory_20_scale_5_imag_tb),
.memory_21_scale_5_imag(memory_21_scale_5_imag_tb),
.memory_22_scale_5_imag(memory_22_scale_5_imag_tb),
.memory_23_scale_5_imag(memory_23_scale_5_imag_tb),
.memory_24_scale_5_imag(memory_24_scale_5_imag_tb),
.memory_25_scale_5_imag(memory_25_scale_5_imag_tb),
.memory_26_scale_5_imag(memory_26_scale_5_imag_tb),
.memory_27_scale_5_imag(memory_27_scale_5_imag_tb),
.memory_28_scale_5_imag(memory_28_scale_5_imag_tb),
.memory_29_scale_5_imag(memory_29_scale_5_imag_tb),
.memory_30_scale_5_imag(memory_30_scale_5_imag_tb),
.memory_31_scale_5_imag(memory_31_scale_5_imag_tb),
.memory_0_scale_6_imag(memory_0_scale_6_imag_tb),
.memory_1_scale_6_imag(memory_1_scale_6_imag_tb),
.memory_2_scale_6_imag(memory_2_scale_6_imag_tb),
.memory_3_scale_6_imag(memory_3_scale_6_imag_tb),
.memory_4_scale_6_imag(memory_4_scale_6_imag_tb),
.memory_5_scale_6_imag(memory_5_scale_6_imag_tb),
.memory_6_scale_6_imag(memory_6_scale_6_imag_tb),
.memory_7_scale_6_imag(memory_7_scale_6_imag_tb),
.memory_8_scale_6_imag(memory_8_scale_6_imag_tb),
.memory_9_scale_6_imag(memory_9_scale_6_imag_tb),
.memory_10_scale_6_imag(memory_10_scale_6_imag_tb),
.memory_11_scale_6_imag(memory_11_scale_6_imag_tb),
.memory_12_scale_6_imag(memory_12_scale_6_imag_tb),
.memory_13_scale_6_imag(memory_13_scale_6_imag_tb),
.memory_14_scale_6_imag(memory_14_scale_6_imag_tb),
.memory_15_scale_6_imag(memory_15_scale_6_imag_tb),
.memory_16_scale_6_imag(memory_16_scale_6_imag_tb),
.memory_17_scale_6_imag(memory_17_scale_6_imag_tb),
.memory_18_scale_6_imag(memory_18_scale_6_imag_tb),
.memory_19_scale_6_imag(memory_19_scale_6_imag_tb),
.memory_20_scale_6_imag(memory_20_scale_6_imag_tb),
.memory_21_scale_6_imag(memory_21_scale_6_imag_tb),
.memory_22_scale_6_imag(memory_22_scale_6_imag_tb),
.memory_23_scale_6_imag(memory_23_scale_6_imag_tb),
.memory_24_scale_6_imag(memory_24_scale_6_imag_tb),
.memory_25_scale_6_imag(memory_25_scale_6_imag_tb),
.memory_26_scale_6_imag(memory_26_scale_6_imag_tb),
.memory_27_scale_6_imag(memory_27_scale_6_imag_tb),
.memory_28_scale_6_imag(memory_28_scale_6_imag_tb),
.memory_29_scale_6_imag(memory_29_scale_6_imag_tb),
.memory_30_scale_6_imag(memory_30_scale_6_imag_tb),
.memory_31_scale_6_imag(memory_31_scale_6_imag_tb),
.memory_0_scale_7_imag(memory_0_scale_7_imag_tb),
.memory_1_scale_7_imag(memory_1_scale_7_imag_tb),
.memory_2_scale_7_imag(memory_2_scale_7_imag_tb),
.memory_3_scale_7_imag(memory_3_scale_7_imag_tb),
.memory_4_scale_7_imag(memory_4_scale_7_imag_tb),
.memory_5_scale_7_imag(memory_5_scale_7_imag_tb),
.memory_6_scale_7_imag(memory_6_scale_7_imag_tb),
.memory_7_scale_7_imag(memory_7_scale_7_imag_tb),
.memory_8_scale_7_imag(memory_8_scale_7_imag_tb),
.memory_9_scale_7_imag(memory_9_scale_7_imag_tb),
.memory_10_scale_7_imag(memory_10_scale_7_imag_tb),
.memory_11_scale_7_imag(memory_11_scale_7_imag_tb),
.memory_12_scale_7_imag(memory_12_scale_7_imag_tb),
.memory_13_scale_7_imag(memory_13_scale_7_imag_tb),
.memory_14_scale_7_imag(memory_14_scale_7_imag_tb),
.memory_15_scale_7_imag(memory_15_scale_7_imag_tb),
.memory_16_scale_7_imag(memory_16_scale_7_imag_tb),
.memory_17_scale_7_imag(memory_17_scale_7_imag_tb),
.memory_18_scale_7_imag(memory_18_scale_7_imag_tb),
.memory_19_scale_7_imag(memory_19_scale_7_imag_tb),
.memory_20_scale_7_imag(memory_20_scale_7_imag_tb),
.memory_21_scale_7_imag(memory_21_scale_7_imag_tb),
.memory_22_scale_7_imag(memory_22_scale_7_imag_tb),
.memory_23_scale_7_imag(memory_23_scale_7_imag_tb),
.memory_24_scale_7_imag(memory_24_scale_7_imag_tb),
.memory_25_scale_7_imag(memory_25_scale_7_imag_tb),
.memory_26_scale_7_imag(memory_26_scale_7_imag_tb),
.memory_27_scale_7_imag(memory_27_scale_7_imag_tb),
.memory_28_scale_7_imag(memory_28_scale_7_imag_tb),
.memory_29_scale_7_imag(memory_29_scale_7_imag_tb),
.memory_30_scale_7_imag(memory_30_scale_7_imag_tb),
.memory_31_scale_7_imag(memory_31_scale_7_imag_tb),
.memory_0_scale_8_imag(memory_0_scale_8_imag_tb),
.memory_1_scale_8_imag(memory_1_scale_8_imag_tb),
.memory_2_scale_8_imag(memory_2_scale_8_imag_tb),
.memory_3_scale_8_imag(memory_3_scale_8_imag_tb),
.memory_4_scale_8_imag(memory_4_scale_8_imag_tb),
.memory_5_scale_8_imag(memory_5_scale_8_imag_tb),
.memory_6_scale_8_imag(memory_6_scale_8_imag_tb),
.memory_7_scale_8_imag(memory_7_scale_8_imag_tb),
.memory_8_scale_8_imag(memory_8_scale_8_imag_tb),
.memory_9_scale_8_imag(memory_9_scale_8_imag_tb),
.memory_10_scale_8_imag(memory_10_scale_8_imag_tb),
.memory_11_scale_8_imag(memory_11_scale_8_imag_tb),
.memory_12_scale_8_imag(memory_12_scale_8_imag_tb),
.memory_13_scale_8_imag(memory_13_scale_8_imag_tb),
.memory_14_scale_8_imag(memory_14_scale_8_imag_tb),
.memory_15_scale_8_imag(memory_15_scale_8_imag_tb),
.memory_16_scale_8_imag(memory_16_scale_8_imag_tb),
.memory_17_scale_8_imag(memory_17_scale_8_imag_tb),
.memory_18_scale_8_imag(memory_18_scale_8_imag_tb),
.memory_19_scale_8_imag(memory_19_scale_8_imag_tb),
.memory_20_scale_8_imag(memory_20_scale_8_imag_tb),
.memory_21_scale_8_imag(memory_21_scale_8_imag_tb),
.memory_22_scale_8_imag(memory_22_scale_8_imag_tb),
.memory_23_scale_8_imag(memory_23_scale_8_imag_tb),
.memory_24_scale_8_imag(memory_24_scale_8_imag_tb),
.memory_25_scale_8_imag(memory_25_scale_8_imag_tb),
.memory_26_scale_8_imag(memory_26_scale_8_imag_tb),
.memory_27_scale_8_imag(memory_27_scale_8_imag_tb),
.memory_28_scale_8_imag(memory_28_scale_8_imag_tb),
.memory_29_scale_8_imag(memory_29_scale_8_imag_tb),
.memory_30_scale_8_imag(memory_30_scale_8_imag_tb),
.memory_31_scale_8_imag(memory_31_scale_8_imag_tb),
.memory_0_scale_9_imag(memory_0_scale_9_imag_tb),
.memory_1_scale_9_imag(memory_1_scale_9_imag_tb),
.memory_2_scale_9_imag(memory_2_scale_9_imag_tb),
.memory_3_scale_9_imag(memory_3_scale_9_imag_tb),
.memory_4_scale_9_imag(memory_4_scale_9_imag_tb),
.memory_5_scale_9_imag(memory_5_scale_9_imag_tb),
.memory_6_scale_9_imag(memory_6_scale_9_imag_tb),
.memory_7_scale_9_imag(memory_7_scale_9_imag_tb),
.memory_8_scale_9_imag(memory_8_scale_9_imag_tb),
.memory_9_scale_9_imag(memory_9_scale_9_imag_tb),
.memory_10_scale_9_imag(memory_10_scale_9_imag_tb),
.memory_11_scale_9_imag(memory_11_scale_9_imag_tb),
.memory_12_scale_9_imag(memory_12_scale_9_imag_tb),
.memory_13_scale_9_imag(memory_13_scale_9_imag_tb),
.memory_14_scale_9_imag(memory_14_scale_9_imag_tb),
.memory_15_scale_9_imag(memory_15_scale_9_imag_tb),
.memory_16_scale_9_imag(memory_16_scale_9_imag_tb),
.memory_17_scale_9_imag(memory_17_scale_9_imag_tb),
.memory_18_scale_9_imag(memory_18_scale_9_imag_tb),
.memory_19_scale_9_imag(memory_19_scale_9_imag_tb),
.memory_20_scale_9_imag(memory_20_scale_9_imag_tb),
.memory_21_scale_9_imag(memory_21_scale_9_imag_tb),
.memory_22_scale_9_imag(memory_22_scale_9_imag_tb),
.memory_23_scale_9_imag(memory_23_scale_9_imag_tb),
.memory_24_scale_9_imag(memory_24_scale_9_imag_tb),
.memory_25_scale_9_imag(memory_25_scale_9_imag_tb),
.memory_26_scale_9_imag(memory_26_scale_9_imag_tb),
.memory_27_scale_9_imag(memory_27_scale_9_imag_tb),
.memory_28_scale_9_imag(memory_28_scale_9_imag_tb),
.memory_29_scale_9_imag(memory_29_scale_9_imag_tb),
.memory_30_scale_9_imag(memory_30_scale_9_imag_tb),
.memory_31_scale_9_imag(memory_31_scale_9_imag_tb),
.memory_0_scale_10_imag(memory_0_scale_10_imag_tb),
.memory_1_scale_10_imag(memory_1_scale_10_imag_tb),
.memory_2_scale_10_imag(memory_2_scale_10_imag_tb),
.memory_3_scale_10_imag(memory_3_scale_10_imag_tb),
.memory_4_scale_10_imag(memory_4_scale_10_imag_tb),
.memory_5_scale_10_imag(memory_5_scale_10_imag_tb),
.memory_6_scale_10_imag(memory_6_scale_10_imag_tb),
.memory_7_scale_10_imag(memory_7_scale_10_imag_tb),
.memory_8_scale_10_imag(memory_8_scale_10_imag_tb),
.memory_9_scale_10_imag(memory_9_scale_10_imag_tb),
.memory_10_scale_10_imag(memory_10_scale_10_imag_tb),
.memory_11_scale_10_imag(memory_11_scale_10_imag_tb),
.memory_12_scale_10_imag(memory_12_scale_10_imag_tb),
.memory_13_scale_10_imag(memory_13_scale_10_imag_tb),
.memory_14_scale_10_imag(memory_14_scale_10_imag_tb),
.memory_15_scale_10_imag(memory_15_scale_10_imag_tb),
.memory_16_scale_10_imag(memory_16_scale_10_imag_tb),
.memory_17_scale_10_imag(memory_17_scale_10_imag_tb),
.memory_18_scale_10_imag(memory_18_scale_10_imag_tb),
.memory_19_scale_10_imag(memory_19_scale_10_imag_tb),
.memory_20_scale_10_imag(memory_20_scale_10_imag_tb),
.memory_21_scale_10_imag(memory_21_scale_10_imag_tb),
.memory_22_scale_10_imag(memory_22_scale_10_imag_tb),
.memory_23_scale_10_imag(memory_23_scale_10_imag_tb),
.memory_24_scale_10_imag(memory_24_scale_10_imag_tb),
.memory_25_scale_10_imag(memory_25_scale_10_imag_tb),
.memory_26_scale_10_imag(memory_26_scale_10_imag_tb),
.memory_27_scale_10_imag(memory_27_scale_10_imag_tb),
.memory_28_scale_10_imag(memory_28_scale_10_imag_tb),
.memory_29_scale_10_imag(memory_29_scale_10_imag_tb),
.memory_30_scale_10_imag(memory_30_scale_10_imag_tb),
.memory_31_scale_10_imag(memory_31_scale_10_imag_tb),
.memory_0_scale_11_imag(memory_0_scale_11_imag_tb),
.memory_1_scale_11_imag(memory_1_scale_11_imag_tb),
.memory_2_scale_11_imag(memory_2_scale_11_imag_tb),
.memory_3_scale_11_imag(memory_3_scale_11_imag_tb),
.memory_4_scale_11_imag(memory_4_scale_11_imag_tb),
.memory_5_scale_11_imag(memory_5_scale_11_imag_tb),
.memory_6_scale_11_imag(memory_6_scale_11_imag_tb),
.memory_7_scale_11_imag(memory_7_scale_11_imag_tb),
.memory_8_scale_11_imag(memory_8_scale_11_imag_tb),
.memory_9_scale_11_imag(memory_9_scale_11_imag_tb),
.memory_10_scale_11_imag(memory_10_scale_11_imag_tb),
.memory_11_scale_11_imag(memory_11_scale_11_imag_tb),
.memory_12_scale_11_imag(memory_12_scale_11_imag_tb),
.memory_13_scale_11_imag(memory_13_scale_11_imag_tb),
.memory_14_scale_11_imag(memory_14_scale_11_imag_tb),
.memory_15_scale_11_imag(memory_15_scale_11_imag_tb),
.memory_16_scale_11_imag(memory_16_scale_11_imag_tb),
.memory_17_scale_11_imag(memory_17_scale_11_imag_tb),
.memory_18_scale_11_imag(memory_18_scale_11_imag_tb),
.memory_19_scale_11_imag(memory_19_scale_11_imag_tb),
.memory_20_scale_11_imag(memory_20_scale_11_imag_tb),
.memory_21_scale_11_imag(memory_21_scale_11_imag_tb),
.memory_22_scale_11_imag(memory_22_scale_11_imag_tb),
.memory_23_scale_11_imag(memory_23_scale_11_imag_tb),
.memory_24_scale_11_imag(memory_24_scale_11_imag_tb),
.memory_25_scale_11_imag(memory_25_scale_11_imag_tb),
.memory_26_scale_11_imag(memory_26_scale_11_imag_tb),
.memory_27_scale_11_imag(memory_27_scale_11_imag_tb),
.memory_28_scale_11_imag(memory_28_scale_11_imag_tb),
.memory_29_scale_11_imag(memory_29_scale_11_imag_tb),
.memory_30_scale_11_imag(memory_30_scale_11_imag_tb),
.memory_31_scale_11_imag(memory_31_scale_11_imag_tb),
.memory_0_scale_12_imag(memory_0_scale_12_imag_tb),
.memory_1_scale_12_imag(memory_1_scale_12_imag_tb),
.memory_2_scale_12_imag(memory_2_scale_12_imag_tb),
.memory_3_scale_12_imag(memory_3_scale_12_imag_tb),
.memory_4_scale_12_imag(memory_4_scale_12_imag_tb),
.memory_5_scale_12_imag(memory_5_scale_12_imag_tb),
.memory_6_scale_12_imag(memory_6_scale_12_imag_tb),
.memory_7_scale_12_imag(memory_7_scale_12_imag_tb),
.memory_8_scale_12_imag(memory_8_scale_12_imag_tb),
.memory_9_scale_12_imag(memory_9_scale_12_imag_tb),
.memory_10_scale_12_imag(memory_10_scale_12_imag_tb),
.memory_11_scale_12_imag(memory_11_scale_12_imag_tb),
.memory_12_scale_12_imag(memory_12_scale_12_imag_tb),
.memory_13_scale_12_imag(memory_13_scale_12_imag_tb),
.memory_14_scale_12_imag(memory_14_scale_12_imag_tb),
.memory_15_scale_12_imag(memory_15_scale_12_imag_tb),
.memory_16_scale_12_imag(memory_16_scale_12_imag_tb),
.memory_17_scale_12_imag(memory_17_scale_12_imag_tb),
.memory_18_scale_12_imag(memory_18_scale_12_imag_tb),
.memory_19_scale_12_imag(memory_19_scale_12_imag_tb),
.memory_20_scale_12_imag(memory_20_scale_12_imag_tb),
.memory_21_scale_12_imag(memory_21_scale_12_imag_tb),
.memory_22_scale_12_imag(memory_22_scale_12_imag_tb),
.memory_23_scale_12_imag(memory_23_scale_12_imag_tb),
.memory_24_scale_12_imag(memory_24_scale_12_imag_tb),
.memory_25_scale_12_imag(memory_25_scale_12_imag_tb),
.memory_26_scale_12_imag(memory_26_scale_12_imag_tb),
.memory_27_scale_12_imag(memory_27_scale_12_imag_tb),
.memory_28_scale_12_imag(memory_28_scale_12_imag_tb),
.memory_29_scale_12_imag(memory_29_scale_12_imag_tb),
.memory_30_scale_12_imag(memory_30_scale_12_imag_tb),
.memory_31_scale_12_imag(memory_31_scale_12_imag_tb),
.memory_0_scale_13_imag(memory_0_scale_13_imag_tb),
.memory_1_scale_13_imag(memory_1_scale_13_imag_tb),
.memory_2_scale_13_imag(memory_2_scale_13_imag_tb),
.memory_3_scale_13_imag(memory_3_scale_13_imag_tb),
.memory_4_scale_13_imag(memory_4_scale_13_imag_tb),
.memory_5_scale_13_imag(memory_5_scale_13_imag_tb),
.memory_6_scale_13_imag(memory_6_scale_13_imag_tb),
.memory_7_scale_13_imag(memory_7_scale_13_imag_tb),
.memory_8_scale_13_imag(memory_8_scale_13_imag_tb),
.memory_9_scale_13_imag(memory_9_scale_13_imag_tb),
.memory_10_scale_13_imag(memory_10_scale_13_imag_tb),
.memory_11_scale_13_imag(memory_11_scale_13_imag_tb),
.memory_12_scale_13_imag(memory_12_scale_13_imag_tb),
.memory_13_scale_13_imag(memory_13_scale_13_imag_tb),
.memory_14_scale_13_imag(memory_14_scale_13_imag_tb),
.memory_15_scale_13_imag(memory_15_scale_13_imag_tb),
.memory_16_scale_13_imag(memory_16_scale_13_imag_tb),
.memory_17_scale_13_imag(memory_17_scale_13_imag_tb),
.memory_18_scale_13_imag(memory_18_scale_13_imag_tb),
.memory_19_scale_13_imag(memory_19_scale_13_imag_tb),
.memory_20_scale_13_imag(memory_20_scale_13_imag_tb),
.memory_21_scale_13_imag(memory_21_scale_13_imag_tb),
.memory_22_scale_13_imag(memory_22_scale_13_imag_tb),
.memory_23_scale_13_imag(memory_23_scale_13_imag_tb),
.memory_24_scale_13_imag(memory_24_scale_13_imag_tb),
.memory_25_scale_13_imag(memory_25_scale_13_imag_tb),
.memory_26_scale_13_imag(memory_26_scale_13_imag_tb),
.memory_27_scale_13_imag(memory_27_scale_13_imag_tb),
.memory_28_scale_13_imag(memory_28_scale_13_imag_tb),
.memory_29_scale_13_imag(memory_29_scale_13_imag_tb),
.memory_30_scale_13_imag(memory_30_scale_13_imag_tb),
.memory_31_scale_13_imag(memory_31_scale_13_imag_tb),
.memory_0_scale_14_imag(memory_0_scale_14_imag_tb),
.memory_1_scale_14_imag(memory_1_scale_14_imag_tb),
.memory_2_scale_14_imag(memory_2_scale_14_imag_tb),
.memory_3_scale_14_imag(memory_3_scale_14_imag_tb),
.memory_4_scale_14_imag(memory_4_scale_14_imag_tb),
.memory_5_scale_14_imag(memory_5_scale_14_imag_tb),
.memory_6_scale_14_imag(memory_6_scale_14_imag_tb),
.memory_7_scale_14_imag(memory_7_scale_14_imag_tb),
.memory_8_scale_14_imag(memory_8_scale_14_imag_tb),
.memory_9_scale_14_imag(memory_9_scale_14_imag_tb),
.memory_10_scale_14_imag(memory_10_scale_14_imag_tb),
.memory_11_scale_14_imag(memory_11_scale_14_imag_tb),
.memory_12_scale_14_imag(memory_12_scale_14_imag_tb),
.memory_13_scale_14_imag(memory_13_scale_14_imag_tb),
.memory_14_scale_14_imag(memory_14_scale_14_imag_tb),
.memory_15_scale_14_imag(memory_15_scale_14_imag_tb),
.memory_16_scale_14_imag(memory_16_scale_14_imag_tb),
.memory_17_scale_14_imag(memory_17_scale_14_imag_tb),
.memory_18_scale_14_imag(memory_18_scale_14_imag_tb),
.memory_19_scale_14_imag(memory_19_scale_14_imag_tb),
.memory_20_scale_14_imag(memory_20_scale_14_imag_tb),
.memory_21_scale_14_imag(memory_21_scale_14_imag_tb),
.memory_22_scale_14_imag(memory_22_scale_14_imag_tb),
.memory_23_scale_14_imag(memory_23_scale_14_imag_tb),
.memory_24_scale_14_imag(memory_24_scale_14_imag_tb),
.memory_25_scale_14_imag(memory_25_scale_14_imag_tb),
.memory_26_scale_14_imag(memory_26_scale_14_imag_tb),
.memory_27_scale_14_imag(memory_27_scale_14_imag_tb),
.memory_28_scale_14_imag(memory_28_scale_14_imag_tb),
.memory_29_scale_14_imag(memory_29_scale_14_imag_tb),
.memory_30_scale_14_imag(memory_30_scale_14_imag_tb),
.memory_31_scale_14_imag(memory_31_scale_14_imag_tb),
.memory_0_scale_15_imag(memory_0_scale_15_imag_tb),
.memory_1_scale_15_imag(memory_1_scale_15_imag_tb),
.memory_2_scale_15_imag(memory_2_scale_15_imag_tb),
.memory_3_scale_15_imag(memory_3_scale_15_imag_tb),
.memory_4_scale_15_imag(memory_4_scale_15_imag_tb),
.memory_5_scale_15_imag(memory_5_scale_15_imag_tb),
.memory_6_scale_15_imag(memory_6_scale_15_imag_tb),
.memory_7_scale_15_imag(memory_7_scale_15_imag_tb),
.memory_8_scale_15_imag(memory_8_scale_15_imag_tb),
.memory_9_scale_15_imag(memory_9_scale_15_imag_tb),
.memory_10_scale_15_imag(memory_10_scale_15_imag_tb),
.memory_11_scale_15_imag(memory_11_scale_15_imag_tb),
.memory_12_scale_15_imag(memory_12_scale_15_imag_tb),
.memory_13_scale_15_imag(memory_13_scale_15_imag_tb),
.memory_14_scale_15_imag(memory_14_scale_15_imag_tb),
.memory_15_scale_15_imag(memory_15_scale_15_imag_tb),
.memory_16_scale_15_imag(memory_16_scale_15_imag_tb),
.memory_17_scale_15_imag(memory_17_scale_15_imag_tb),
.memory_18_scale_15_imag(memory_18_scale_15_imag_tb),
.memory_19_scale_15_imag(memory_19_scale_15_imag_tb),
.memory_20_scale_15_imag(memory_20_scale_15_imag_tb),
.memory_21_scale_15_imag(memory_21_scale_15_imag_tb),
.memory_22_scale_15_imag(memory_22_scale_15_imag_tb),
.memory_23_scale_15_imag(memory_23_scale_15_imag_tb),
.memory_24_scale_15_imag(memory_24_scale_15_imag_tb),
.memory_25_scale_15_imag(memory_25_scale_15_imag_tb),
.memory_26_scale_15_imag(memory_26_scale_15_imag_tb),
.memory_27_scale_15_imag(memory_27_scale_15_imag_tb),
.memory_28_scale_15_imag(memory_28_scale_15_imag_tb),
.memory_29_scale_15_imag(memory_29_scale_15_imag_tb),
.memory_30_scale_15_imag(memory_30_scale_15_imag_tb),
.memory_31_scale_15_imag(memory_31_scale_15_imag_tb)


);


	always #(Clock_Period / 2) clk_tb = ~clk_tb ;
	
	initial begin
	$dumpfile("CWT.vcd");
	$dumpvars;

  reset();
	initialize();
	
  
	/* TEST CASE 1 */
	//TEST_CASE_1();
	
	TEST_CASE_2();
  FFT_Operation();

	#(10 * Clock_Period)
	$stop ;

end


task initialize ;
begin
  ready_inputs_tb = 1'b0;
  clk_tb = 1'b1 ; 
  rst_tb = 1'b1;
  read_scale_ram_addresses = 2'b00;
x0_r_tb = 16'b00000000_00000000;
x0_i_tb = 16'b00000000_00000000;
x1_r_tb = 16'b00000000_00000000;
x1_i_tb = 16'b00000000_00000000;
x2_r_tb = 16'b00000000_00000000;
x2_i_tb = 16'b00000000_00000000;
x3_r_tb = 16'b00000000_00000000;
x3_i_tb = 16'b00000000_00000000;
x4_r_tb = 16'b00000000_00000000;
x4_i_tb = 16'b00000000_00000000;
x5_r_tb = 16'b00000000_00000000;
x5_i_tb = 16'b00000000_00000000;
x6_r_tb = 16'b00000000_00000000;
x6_i_tb = 16'b00000000_00000000;
x7_r_tb = 16'b00000000_00000000;
x7_i_tb = 16'b00000000_00000000;
x8_r_tb = 16'b00000000_00000000;
x8_i_tb = 16'b00000000_00000000;
x9_r_tb = 16'b00000000_00000000;
x9_i_tb = 16'b00000000_00000000;
x10_r_tb = 16'b00000000_00000000;
x10_i_tb = 16'b00000000_00000000;
x11_r_tb = 16'b00000000_00000000;
x11_i_tb = 16'b00000000_00000000;
x12_r_tb = 16'b00000000_00000000;
x12_i_tb = 16'b00000000_00000000;
x13_r_tb = 16'b00000000_00000000;
x13_i_tb = 16'b00000000_00000000;
x14_r_tb = 16'b00000000_00000000;
x14_i_tb = 16'b00000000_00000000;
x15_r_tb = 16'b00000000_00000000;
x15_i_tb = 16'b00000000_00000000;
x16_r_tb = 16'b00000000_00000000;
x16_i_tb = 16'b00000000_00000000;
x17_r_tb = 16'b00000000_00000000;
x17_i_tb = 16'b00000000_00000000;
x18_r_tb = 16'b00000000_00000000;
x18_i_tb = 16'b00000000_00000000;
x19_r_tb = 16'b00000000_00000000;
x19_i_tb = 16'b00000000_00000000;
x20_r_tb = 16'b00000000_00000000;
x20_i_tb = 16'b00000000_00000000;
x21_r_tb = 16'b00000000_00000000;
x21_i_tb = 16'b00000000_00000000;
x22_r_tb = 16'b00000000_00000000;
x22_i_tb = 16'b00000000_00000000;
x23_r_tb = 16'b00000000_00000000;
x23_i_tb = 16'b00000000_00000000;
x24_r_tb = 16'b00000000_00000000;
x24_i_tb = 16'b00000000_00000000;
x25_r_tb = 16'b00000000_00000000;
x25_i_tb = 16'b00000000_00000000;
x26_r_tb = 16'b00000000_00000000;
x26_i_tb = 16'b00000000_00000000;
x27_r_tb = 16'b00000000_00000000;
x27_i_tb = 16'b00000000_00000000;
x28_r_tb = 16'b00000000_00000000;
x28_i_tb = 16'b00000000_00000000;
x29_r_tb = 16'b00000000_00000000;
x29_i_tb = 16'b00000000_00000000;
x30_r_tb = 16'b00000000_00000000;
x30_i_tb = 16'b00000000_00000000;
x31_r_tb = 16'b00000000_00000000;
x31_i_tb = 16'b00000000_00000000;
x32_r_tb = 16'b00000000_00000000;
x32_i_tb = 16'b00000000_00000000;
x33_r_tb = 16'b00000000_00000000;
x33_i_tb = 16'b00000000_00000000;
x34_r_tb = 16'b00000000_00000000;
x34_i_tb = 16'b00000000_00000000;
x35_r_tb = 16'b00000000_00000000;
x35_i_tb = 16'b00000000_00000000;
x36_r_tb = 16'b00000000_00000000;
x36_i_tb = 16'b00000000_00000000;
x37_r_tb = 16'b00000000_00000000;
x37_i_tb = 16'b00000000_00000000;
x38_r_tb = 16'b00000000_00000000;
x38_i_tb = 16'b00000000_00000000;
x39_r_tb = 16'b00000000_00000000;
x39_i_tb = 16'b00000000_00000000;
x40_r_tb = 16'b00000000_00000000;
x40_i_tb = 16'b00000000_00000000;
x41_r_tb = 16'b00000000_00000000;
x41_i_tb = 16'b00000000_00000000;
x42_r_tb = 16'b00000000_00000000;
x42_i_tb = 16'b00000000_00000000;
x43_r_tb = 16'b00000000_00000000;
x43_i_tb = 16'b00000000_00000000;
x44_r_tb = 16'b00000000_00000000;
x44_i_tb = 16'b00000000_00000000;
x45_r_tb = 16'b00000000_00000000;
x45_i_tb = 16'b00000000_00000000;
x46_r_tb = 16'b00000000_00000000;
x46_i_tb = 16'b00000000_00000000;
x47_r_tb = 16'b00000000_00000000;
x47_i_tb = 16'b00000000_00000000;
x48_r_tb = 16'b00000000_00000000;
x48_i_tb = 16'b00000000_00000000;
x49_r_tb = 16'b00000000_00000000;
x49_i_tb = 16'b00000000_00000000;
x50_r_tb = 16'b00000000_00000000;
x50_i_tb = 16'b00000000_00000000;
x51_r_tb = 16'b00000000_00000000;
x51_i_tb = 16'b00000000_00000000;
x52_r_tb = 16'b00000000_00000000;
x52_i_tb = 16'b00000000_00000000;
x53_r_tb = 16'b00000000_00000000;
x53_i_tb = 16'b00000000_00000000;
x54_r_tb = 16'b00000000_00000000;
x54_i_tb = 16'b00000000_00000000;
x55_r_tb = 16'b00000000_00000000;
x55_i_tb = 16'b00000000_00000000;
x56_r_tb = 16'b00000000_00000000;
x56_i_tb = 16'b00000000_00000000;
x57_r_tb = 16'b00000000_00000000;
x57_i_tb = 16'b00000000_00000000;
x58_r_tb = 16'b00000000_00000000;
x58_i_tb = 16'b00000000_00000000;
x59_r_tb = 16'b00000000_00000000;
x59_i_tb = 16'b00000000_00000000;
x60_r_tb = 16'b00000000_00000000;
x60_i_tb = 16'b00000000_00000000;
x61_r_tb = 16'b00000000_00000000;
x61_i_tb = 16'b00000000_00000000;
x62_r_tb = 16'b00000000_00000000;
x62_i_tb = 16'b00000000_00000000;
x63_r_tb = 16'b00000000_00000000;
x63_i_tb = 16'b00000000_00000000;
x64_r_tb = 16'b00000000_00000000;
x64_i_tb = 16'b00000000_00000000;
x65_r_tb = 16'b00000000_00000000;
x65_i_tb = 16'b00000000_00000000;
x66_r_tb = 16'b00000000_00000000;
x66_i_tb = 16'b00000000_00000000;
x67_r_tb = 16'b00000000_00000000;
x67_i_tb = 16'b00000000_00000000;
x68_r_tb = 16'b00000000_00000000;
x68_i_tb = 16'b00000000_00000000;
x69_r_tb = 16'b00000000_00000000;
x69_i_tb = 16'b00000000_00000000;
x70_r_tb = 16'b00000000_00000000;
x70_i_tb = 16'b00000000_00000000;
x71_r_tb = 16'b00000000_00000000;
x71_i_tb = 16'b00000000_00000000;
x72_r_tb = 16'b00000000_00000000;
x72_i_tb = 16'b00000000_00000000;
x73_r_tb = 16'b00000000_00000000;
x73_i_tb = 16'b00000000_00000000;
x74_r_tb = 16'b00000000_00000000;
x74_i_tb = 16'b00000000_00000000;
x75_r_tb = 16'b00000000_00000000;
x75_i_tb = 16'b00000000_00000000;
x76_r_tb = 16'b00000000_00000000;
x76_i_tb = 16'b00000000_00000000;
x77_r_tb = 16'b00000000_00000000;
x77_i_tb = 16'b00000000_00000000;
x78_r_tb = 16'b00000000_00000000;
x78_i_tb = 16'b00000000_00000000;
x79_r_tb = 16'b00000000_00000000;
x79_i_tb = 16'b00000000_00000000;
x80_r_tb = 16'b00000000_00000000;
x80_i_tb = 16'b00000000_00000000;
x81_r_tb = 16'b00000000_00000000;
x81_i_tb = 16'b00000000_00000000;
x82_r_tb = 16'b00000000_00000000;
x82_i_tb = 16'b00000000_00000000;
x83_r_tb = 16'b00000000_00000000;
x83_i_tb = 16'b00000000_00000000;
x84_r_tb = 16'b00000000_00000000;
x84_i_tb = 16'b00000000_00000000;
x85_r_tb = 16'b00000000_00000000;
x85_i_tb = 16'b00000000_00000000;
x86_r_tb = 16'b00000000_00000000;
x86_i_tb = 16'b00000000_00000000;
x87_r_tb = 16'b00000000_00000000;
x87_i_tb = 16'b00000000_00000000;
x88_r_tb = 16'b00000000_00000000;
x88_i_tb = 16'b00000000_00000000;
x89_r_tb = 16'b00000000_00000000;
x89_i_tb = 16'b00000000_00000000;
x90_r_tb = 16'b00000000_00000000;
x90_i_tb = 16'b00000000_00000000;
x91_r_tb = 16'b00000000_00000000;
x91_i_tb = 16'b00000000_00000000;
x92_r_tb = 16'b00000000_00000000;
x92_i_tb = 16'b00000000_00000000;
x93_r_tb = 16'b00000000_00000000;
x93_i_tb = 16'b00000000_00000000;
x94_r_tb = 16'b00000000_00000000;
x94_i_tb = 16'b00000000_00000000;
x95_r_tb = 16'b00000000_00000000;
x95_i_tb = 16'b00000000_00000000;
x96_r_tb = 16'b00000000_00000000;
x96_i_tb = 16'b00000000_00000000;
x97_r_tb = 16'b00000000_00000000;
x97_i_tb = 16'b00000000_00000000;
x98_r_tb = 16'b00000000_00000000;
x98_i_tb = 16'b00000000_00000000;
x99_r_tb = 16'b00000000_00000000;
x99_i_tb = 16'b00000000_00000000;
x100_r_tb = 16'b00000000_00000000;
x100_i_tb = 16'b00000000_00000000;
x101_r_tb = 16'b00000000_00000000;
x101_i_tb = 16'b00000000_00000000;
x102_r_tb = 16'b00000000_00000000;
x102_i_tb = 16'b00000000_00000000;
x103_r_tb = 16'b00000000_00000000;
x103_i_tb = 16'b00000000_00000000;
x104_r_tb = 16'b00000000_00000000;
x104_i_tb = 16'b00000000_00000000;
x105_r_tb = 16'b00000000_00000000;
x105_i_tb = 16'b00000000_00000000;
x106_r_tb = 16'b00000000_00000000;
x106_i_tb = 16'b00000000_00000000;
x107_r_tb = 16'b00000000_00000000;
x107_i_tb = 16'b00000000_00000000;
x108_r_tb = 16'b00000000_00000000;
x108_i_tb = 16'b00000000_00000000;
x109_r_tb = 16'b00000000_00000000;
x109_i_tb = 16'b00000000_00000000;
x110_r_tb = 16'b00000000_00000000;
x110_i_tb = 16'b00000000_00000000;
x111_r_tb = 16'b00000000_00000000;
x111_i_tb = 16'b00000000_00000000;
x112_r_tb = 16'b00000000_00000000;
x112_i_tb = 16'b00000000_00000000;
x113_r_tb = 16'b00000000_00000000;
x113_i_tb = 16'b00000000_00000000;
x114_r_tb = 16'b00000000_00000000;
x114_i_tb = 16'b00000000_00000000;
x115_r_tb = 16'b00000000_00000000;
x115_i_tb = 16'b00000000_00000000;
x116_r_tb = 16'b00000000_00000000;
x116_i_tb = 16'b00000000_00000000;
x117_r_tb = 16'b00000000_00000000;
x117_i_tb = 16'b00000000_00000000;
x118_r_tb = 16'b00000000_00000000;
x118_i_tb = 16'b00000000_00000000;
x119_r_tb = 16'b00000000_00000000;
x119_i_tb = 16'b00000000_00000000;
x120_r_tb = 16'b00000000_00000000;
x120_i_tb = 16'b00000000_00000000;
x121_r_tb = 16'b00000000_00000000;
x121_i_tb = 16'b00000000_00000000;
x122_r_tb = 16'b00000000_00000000;
x122_i_tb = 16'b00000000_00000000;
x123_r_tb = 16'b00000000_00000000;
x123_i_tb = 16'b00000000_00000000;
x124_r_tb = 16'b00000000_00000000;
x124_i_tb = 16'b00000000_00000000;
x125_r_tb = 16'b00000000_00000000;
x125_i_tb = 16'b00000000_00000000;
x126_r_tb = 16'b00000000_00000000;
x126_i_tb = 16'b00000000_00000000;
x127_r_tb = 16'b00000000_00000000;
x127_i_tb = 16'b00000000_00000000;
end
endtask

task reset ;
  begin
	/* Reset */
    #(Clock_Period)
    rst_tb = 1'b0 ;
    #(Clock_Period)
    rst_tb = 1'b1 ;
  end
endtask



task TEST_CASE_1;
  begin
	/* TEST CASE 2 */
  x0_r_tb = 16'b11111111_11011011;
x0_i_tb =16'b11111111_11110000;
x1_r_tb = 16'b11111111_11011011;
x1_i_tb =16'b11111111_11110000;
x2_r_tb = 16'b11111111_11011011;
x2_i_tb =16'b11111111_11110000;
x3_r_tb = 16'b11111111_11011011;
x3_i_tb =16'b11111111_11110000;
x4_r_tb = 16'b11111111_11011011;
x4_i_tb =16'b11111111_11110000;
x5_r_tb = 16'b11111111_11011011;
x5_i_tb =16'b11111111_11110000;
x6_r_tb = 16'b11111111_11011011;
x6_i_tb =16'b11111111_11110000;
x7_r_tb = 16'b11111111_11011011;
x7_i_tb =16'b11111111_11110000;
x8_r_tb = 16'b11111111_11011011;
x8_i_tb =16'b11111111_11110000;
    x9_r_tb = 16'b11111111_11100010;
   x9_i_tb = 16'b00000000_00010100;
   x10_r_tb = 16'b00000000_00100010;
   x10_i_tb = 16'b00000000_00010100;
   x11_r_tb = 16'b11111111_11011011;
   x11_i_tb = 16'b11111111_11101011;
   x12_r_tb = 16'b00000000_00100110;
   x12_i_tb = 16'b11111111_11101011;
   x13_r_tb = 16'b11111111_11011000;
   x13_i_tb = 16'b00000000_00010011;
   x14_r_tb = 16'b00000000_00100111;
   x14_i_tb = 16'b00000000_00010001;
   x15_r_tb = 16'b00000000_00101000;
   x15_i_tb = 16'b00000000_00010001;
   x16_r_tb = 16'b11111111_11010100;
   x16_i_tb = 16'b11111111_11110000;
   x17_r_tb = 16'b00000000_00101110;
   x17_i_tb = 16'b11111111_11110010;
   x18_r_tb = 16'b11111111_11010001;
   x18_i_tb = 16'b00000000_00001100;
   x19_r_tb = 16'b00000000_00101011;
   x19_i_tb = 16'b00000000_00001100;
   x20_r_tb = 16'b00000000_00100111;
   x20_i_tb = 16'b00000000_00001010;
   x21_r_tb = 16'b11111111_11010100;
   x21_i_tb = 16'b00000000_00001010;
   x22_r_tb = 16'b11111111_11010010;
   x22_i_tb = 16'b11111111_11110010;
   x23_r_tb = 16'b00000000_00110000;
   x23_i_tb = 16'b11111111_11101101;
   x24_r_tb = 16'b11111111_11010010;
   x24_i_tb = 16'b00000000_00010100;
   x25_r_tb = 16'b00000000_00100111;
   x25_i_tb = 16'b11111111_11101011;
   x26_r_tb = 16'b00000000_00100010;
   x26_i_tb = 16'b00000000_00010001;
   x27_r_tb = 16'b00000000_00100111;
   x27_i_tb = 16'b00000000_00010100;
   x28_r_tb = 16'b00000000_00110000;
   x28_i_tb = 16'b11111111_11101100;
   x29_r_tb = 16'b11111111_11001100;
   x29_i_tb = 16'b00000000_00010111;
   x30_r_tb = 16'b00000000_00111100;
   x30_i_tb = 16'b00000000_00011000;
   x31_r_tb = 16'b11111111_11000111;
   x31_i_tb = 16'b00000000_00010111; 
    x32_r_tb = 16'b11111111_11011011;
x32_i_tb =16'b11111111_11110000;
x33_r_tb = 16'b11111111_11011011;
x33_i_tb =16'b11111111_11110000;
x34_r_tb = 16'b11111111_11011011;
x34_i_tb =16'b11111111_11110000;
x35_r_tb = 16'b11111111_11011011;
x35_i_tb =16'b11111111_11110000;
x36_r_tb = 16'b11111111_11011011;
x36_i_tb =16'b11111111_11110000;
x37_r_tb = 16'b11111111_11011011;
x37_i_tb =16'b11111111_11110000;
x38_r_tb = 16'b11111111_11011011;
x38_i_tb =16'b11111111_11110000;
x39_r_tb = 16'b11111111_11011011;
x39_i_tb =16'b11111111_11110000;
x40_r_tb = 16'b11111111_11011011;
x40_i_tb =16'b11111111_11110000;
    x41_r_tb = 16'b11111111_11100010;
   x41_i_tb = 16'b00000000_00010100;
   x42_r_tb = 16'b00000000_00100010;
   x42_i_tb = 16'b00000000_00010100;
   x43_r_tb = 16'b11111111_11011011;
   x43_i_tb = 16'b11111111_11101011;
   x44_r_tb = 16'b00000000_00100110;
   x44_i_tb = 16'b11111111_11101011;
   x45_r_tb = 16'b11111111_11011000;
   x45_i_tb = 16'b00000000_00010011;
   x46_r_tb = 16'b00000000_00100111;
   x46_i_tb = 16'b00000000_00010001;
   x47_r_tb = 16'b00000000_00101000;
   x47_i_tb = 16'b00000000_00010001;
   x48_r_tb = 16'b11111111_11010100;
   x48_i_tb = 16'b11111111_11110000;
   x49_r_tb = 16'b00000000_00101110;
   x49_i_tb = 16'b11111111_11110010;
   x50_r_tb = 16'b11111111_11010001;
   x50_i_tb = 16'b00000000_00001100;
   x51_r_tb = 16'b00000000_00101011;
   x51_i_tb = 16'b00000000_00001100;
   x52_r_tb = 16'b00000000_00100111;
   x52_i_tb = 16'b00000000_00001010;
   x53_r_tb = 16'b11111111_11010100;
   x53_i_tb = 16'b00000000_00001010;
   x54_r_tb = 16'b11111111_11010010;
   x54_i_tb = 16'b11111111_11110010;
   x55_r_tb = 16'b00000000_00110000;
   x55_i_tb = 16'b11111111_11101101;
   x56_r_tb = 16'b11111111_11010010;
   x56_i_tb = 16'b00000000_00010100;
   x57_r_tb = 16'b00000000_00100111;
   x57_i_tb = 16'b11111111_11101011;
   x58_r_tb = 16'b00000000_00100010;
   x58_i_tb = 16'b00000000_00010001;
   x59_r_tb = 16'b00000000_00100111;
   x59_i_tb = 16'b00000000_00010100;
   x60_r_tb = 16'b00000000_00110000;
   x60_i_tb = 16'b11111111_11101100;
   x61_r_tb = 16'b11111111_11001100;
   x61_i_tb = 16'b00000000_00010111;
   x62_r_tb = 16'b00000000_00111100;
   x62_i_tb = 16'b00000000_00011000;
   x63_r_tb = 16'b11111111_11000111;
   x63_i_tb = 16'b00000000_00010111; 
    x64_r_tb = 16'b11111111_11011011;
x64_i_tb =16'b11111111_11110000;
x65_r_tb = 16'b11111111_11011011;
x65_i_tb =16'b11111111_11110000;
x66_r_tb = 16'b11111111_11011011;
x66_i_tb =16'b11111111_11110000;
x67_r_tb = 16'b11111111_11011011;
x67_i_tb =16'b11111111_11110000;
x68_r_tb = 16'b11111111_11011011;
x68_i_tb =16'b11111111_11110000;
x69_r_tb = 16'b11111111_11011011;
x69_i_tb =16'b11111111_11110000;
x70_r_tb = 16'b11111111_11011011;
x70_i_tb =16'b11111111_11110000;
x71_r_tb = 16'b11111111_11011011;
x71_i_tb =16'b11111111_11110000;
x72_r_tb = 16'b11111111_11011011;
x72_i_tb =16'b11111111_11110000;
    x73_r_tb = 16'b11111111_11100010;
   x73_i_tb = 16'b00000000_00010100;
   x74_r_tb = 16'b00000000_00100010;
   x74_i_tb = 16'b00000000_00010100;
   x75_r_tb = 16'b11111111_11011011;
   x75_i_tb = 16'b11111111_11101011;
   x76_r_tb = 16'b00000000_00100110;
   x76_i_tb = 16'b11111111_11101011;
   x77_r_tb = 16'b11111111_11011000;
   x77_i_tb = 16'b00000000_00010011;
   x78_r_tb = 16'b00000000_00100111;
   x78_i_tb = 16'b00000000_00010001;
   x79_r_tb = 16'b00000000_00101000;
   x79_i_tb = 16'b00000000_00010001;
   x80_r_tb = 16'b11111111_11010100;
   x80_i_tb = 16'b11111111_11110000;
   x81_r_tb = 16'b00000000_00101110;
   x81_i_tb = 16'b11111111_11110010;
   x82_r_tb = 16'b11111111_11010001;
   x82_i_tb = 16'b00000000_00001100;
   x83_r_tb = 16'b00000000_00101011;
   x83_i_tb = 16'b00000000_00001100;
   x84_r_tb = 16'b00000000_00100111;
   x84_i_tb = 16'b00000000_00001010;
   x85_r_tb = 16'b11111111_11010100;
   x85_i_tb = 16'b00000000_00001010;
   x86_r_tb = 16'b11111111_11010010;
   x86_i_tb = 16'b11111111_11110010;
   x87_r_tb = 16'b00000000_00110000;
   x87_i_tb = 16'b11111111_11101101;
   x88_r_tb = 16'b11111111_11010010;
   x88_i_tb = 16'b00000000_00010100;
   x89_r_tb = 16'b00000000_00100111;
   x89_i_tb = 16'b11111111_11101011;
   x90_r_tb = 16'b00000000_00100010;
   x90_i_tb = 16'b00000000_00010001;
   x91_r_tb = 16'b00000000_00100111;
   x91_i_tb = 16'b00000000_00010100;
   x92_r_tb = 16'b00000000_00110000;
   x92_i_tb = 16'b11111111_11101100;
   x93_r_tb = 16'b11111111_11001100;
   x93_i_tb = 16'b00000000_00010111;
   x94_r_tb = 16'b00000000_00111100;
   x94_i_tb = 16'b00000000_00011000;
   x95_r_tb = 16'b11111111_11000111;
   x95_i_tb = 16'b00000000_00010111; 
    x96_r_tb = 16'b11111111_11011011;
x96_i_tb =16'b11111111_11110000;
x97_r_tb = 16'b11111111_11011011;
x97_i_tb =16'b11111111_11110000;
x98_r_tb = 16'b11111111_11011011;
x98_i_tb =16'b11111111_11110000;
x99_r_tb = 16'b11111111_11011011;
x99_i_tb =16'b11111111_11110000;
x100_r_tb = 16'b11111111_11011011;
x100_i_tb =16'b11111111_11110000;
x101_r_tb = 16'b11111111_11011011;
x101_i_tb =16'b11111111_11110000;
x102_r_tb = 16'b11111111_11011011;
x102_i_tb =16'b11111111_11110000;
x103_r_tb = 16'b11111111_11011011;
x103_i_tb =16'b11111111_11110000;
x104_r_tb = 16'b11111111_11011011;
x104_i_tb =16'b11111111_11110000;
    x105_r_tb = 16'b11111111_11100010;
   x105_i_tb = 16'b00000000_00010100;
   x106_r_tb = 16'b00000000_00100010;
   x106_i_tb = 16'b00000000_00010100;
   x107_r_tb = 16'b11111111_11011011;
   x107_i_tb = 16'b11111111_11101011;
   x108_r_tb = 16'b00000000_00100110;
   x108_i_tb = 16'b11111111_11101011;
   x109_r_tb = 16'b11111111_11011000;
   x109_i_tb = 16'b00000000_00010011;
   x110_r_tb = 16'b00000000_00100111;
   x110_i_tb = 16'b00000000_00010001;
   x111_r_tb = 16'b00000000_00101000;
   x111_i_tb = 16'b00000000_00010001;
   x112_r_tb = 16'b11111111_11010100;
   x112_i_tb = 16'b11111111_11110000;
   x113_r_tb = 16'b00000000_00101110;
   x113_i_tb = 16'b11111111_11110010;
   x114_r_tb = 16'b11111111_11010001;
   x114_i_tb = 16'b00000000_00001100;
   x115_r_tb = 16'b00000000_00101011;
   x115_i_tb = 16'b00000000_00001100;
   x116_r_tb = 16'b00000000_00100111;
   x116_i_tb = 16'b00000000_00001010;
   x117_r_tb = 16'b11111111_11010100;
   x117_i_tb = 16'b00000000_00001010;
   x118_r_tb = 16'b11111111_11010010;
   x118_i_tb = 16'b11111111_11110010;
   x119_r_tb = 16'b00000000_00110000;
   x119_i_tb = 16'b11111111_11101101;
   x120_r_tb = 16'b11111111_11010010;
   x120_i_tb = 16'b00000000_00010100;
   x121_r_tb = 16'b00000000_00100111;
   x121_i_tb = 16'b11111111_11101011;
   x122_r_tb = 16'b00000000_00100010;
   x122_i_tb = 16'b00000000_00010001;
   x123_r_tb = 16'b00000000_00100111;
   x123_i_tb = 16'b00000000_00010100;
   x124_r_tb = 16'b00000000_00110000;
   x124_i_tb = 16'b11111111_11101100;
   x125_r_tb = 16'b11111111_11001100;
   x125_i_tb = 16'b00000000_00010111;
   x126_r_tb = 16'b00000000_00111100;
   x126_i_tb = 16'b00000000_00011000;
   x127_r_tb = 16'b11111111_11000111;
   x127_i_tb = 16'b00000000_00010111; 
 
   ready_inputs_tb = 1'b1 ;
    #(4*Clock_Period)
   ready_inputs_tb = 1'b0 ;


  end
endtask

task TEST_CASE_2;
  begin
	/* TEST CASE 2 */
  x0_r_tb = 16'b1111111111011010;
x0_i_tb =16'b0;
x1_r_tb = 16'b1111111111011010;
x1_i_tb =16'b0;
x2_r_tb = 16'b1111111111011010;
x2_i_tb =16'b0;
x3_r_tb = 16'b1111111111011010;
x3_i_tb =16'b0;
x4_r_tb = 16'b1111111111011010;
x4_i_tb =16'b0;
x5_r_tb = 16'b1111111111011010;
x5_i_tb =16'b0;
x6_r_tb = 16'b1111111111011010;
x6_i_tb =16'b0;
x7_r_tb = 16'b1111111111011010;
x7_i_tb =16'b0;
x8_r_tb = 16'b1111111111100001;
x8_i_tb =16'b0;
    x9_r_tb = 16'b1111111111011101;
   x9_i_tb = 16'b0;
   x10_r_tb = 16'b1111111111011010;
   x10_i_tb = 16'b0;
   x11_r_tb = 16'b1111111111011001;
   x11_i_tb = 16'b0;
   x12_r_tb = 16'b1111111111010111;
   x12_i_tb = 16'b0;
   x13_r_tb = 16'b1111111111011000;
   x13_i_tb = 16'b0;
   x14_r_tb = 16'b1111111111010111;
   x14_i_tb = 16'b0;
   x15_r_tb = 16'b1111111111010011;
   x15_i_tb = 16'b0;
   x16_r_tb = 16'b1111111111010001;
   x16_i_tb = 16'b0;
   x17_r_tb = 16'b1111111111010000;
   x17_i_tb = 16'b0;
   x18_r_tb = 16'b1111111111010100;
   x18_i_tb = 16'b0;
   x19_r_tb = 16'b1111111111011000;
   x19_i_tb = 16'b0;
   x20_r_tb = 16'b1111111111010011;
   x20_i_tb = 16'b0;
   x21_r_tb = 16'b1111111111010001;
   x21_i_tb = 16'b0;
   x22_r_tb = 16'b1111111111001111;
   x22_i_tb = 16'b0;
   x23_r_tb = 16'b1111111111010001;
   x23_i_tb = 16'b0;
   x24_r_tb = 16'b1111111111011000;
   x24_i_tb = 16'b0;
   x25_r_tb = 16'b1111111111011101;
   x25_i_tb = 16'b0;
   x26_r_tb = 16'b1111111111011000;
   x26_i_tb = 16'b0;
   x27_r_tb = 16'b1111111111001111;
   x27_i_tb = 16'b0;
   x28_r_tb = 16'b1111111111001011;
   x28_i_tb = 16'b0;
   x29_r_tb = 16'b1111111111000011;
   x29_i_tb = 16'b0;
   x30_r_tb = 16'b1111111111000110;
   x30_i_tb = 16'b0;
   x31_r_tb = 16'b1111111111000001;
   x31_i_tb = 16'b0; 
    x32_r_tb = 16'b1111111111000000;
x32_i_tb =16'b0;
x33_r_tb = 16'b1111111110111101;
x33_i_tb =16'b0;
x34_r_tb = 16'b1111111110111001;
x34_i_tb =16'b0;
x35_r_tb = 16'b1111111110111001;
x35_i_tb =16'b0;
x36_r_tb = 16'b1111111110111001;
x36_i_tb =16'b0;
x37_r_tb = 16'b1111111110111100;
x37_i_tb =16'b0;
x38_r_tb = 16'b1111111110111110;
x38_i_tb =16'b0;
x39_r_tb = 16'b1111111110111100;
x39_i_tb =16'b0;
x40_r_tb = 16'b1111111110111001;
x40_i_tb =16'b0;
    x41_r_tb = 16'b1111111110110101;
   x41_i_tb = 16'b0;
   x42_r_tb = 16'b1111111110110101;
   x42_i_tb = 16'b0;
   x43_r_tb = 16'b1111111110110101;
   x43_i_tb = 16'b0;
   x44_r_tb = 16'b1111111110110101;
   x44_i_tb = 16'b0;
   x45_r_tb = 16'b1111111110110111;
   x45_i_tb = 16'b0;
   x46_r_tb = 16'b1111111110110100;
   x46_i_tb = 16'b0;
   x47_r_tb = 16'b1111111110110001;
   x47_i_tb = 16'b0;
   x48_r_tb = 16'b1111111110110111;
   x48_i_tb = 16'b0;
   x49_r_tb = 16'b1111111110111001;
   x49_i_tb = 16'b0;
   x50_r_tb = 16'b1111111110111001;
   x50_i_tb = 16'b0;
   x51_r_tb = 16'b1111111110111000;
   x51_i_tb = 16'b0;
   x52_r_tb = 16'b1111111110110111;
   x52_i_tb = 16'b0;
   x53_r_tb = 16'b1111111110110001;
   x53_i_tb = 16'b0;
   x54_r_tb = 16'b1111111110110101;
   x54_i_tb = 16'b0;
   x55_r_tb = 16'b1111111110110011;
   x55_i_tb = 16'b0;
   x56_r_tb = 16'b1111111110111000;
   x56_i_tb = 16'b0;
   x57_r_tb = 16'b1111111110110101;
   x57_i_tb = 16'b0;
   x58_r_tb = 16'b1111111110110011;
   x58_i_tb = 16'b0;
   x59_r_tb = 16'b1111111110101111;
   x59_i_tb = 16'b0;
   x60_r_tb = 16'b1111111110101110;
   x60_i_tb = 16'b0;
   x61_r_tb = 16'b1111111110101010;
   x61_i_tb = 16'b0;
   x62_r_tb = 16'b1111111110100011;
   x62_i_tb = 16'b0;
   x63_r_tb = 16'b1111111110011101;
   x63_i_tb = 16'b0; 
    x64_r_tb = 16'b1111111110011101;
x64_i_tb =16'b0;
x65_r_tb = 16'b1111111110011000;
x65_i_tb =16'b0;
x66_r_tb = 16'b1111111110001011;
x66_i_tb =16'b0;
x67_r_tb = 16'b1111111110000011;
x67_i_tb =16'b0;
x68_r_tb = 16'b1111111110000011;
x68_i_tb =16'b0;
x69_r_tb = 16'b1111111110010011;
x69_i_tb =16'b0;
x70_r_tb = 16'b1111111110101011;
x70_i_tb =16'b0;
x71_r_tb = 16'b1111111111000111;
x71_i_tb =16'b0;
x72_r_tb = 16'b1111111111101110;
x72_i_tb =16'b0;
    x73_r_tb = 16'b0000000000011110;
   x73_i_tb = 16'b0;
   x74_r_tb = 16'b0000000001100000;
   x74_i_tb = 16'b0;
   x75_r_tb = 16'b0000000010011110;
   x75_i_tb = 16'b0;
   x76_r_tb = 16'b0000000011000111;
   x76_i_tb = 16'b0;
   x77_r_tb = 16'b0000000011010111;
   x77_i_tb = 16'b0;
   x78_r_tb = 16'b0000000011000011;
   x78_i_tb = 16'b0;
   x79_r_tb = 16'b0000000010000101;
   x79_i_tb = 16'b0;
   x80_r_tb = 16'b0000000000101011;
   x80_i_tb = 16'b0;
   x81_r_tb = 16'b1111111111010101;
   x81_i_tb = 16'b0;
   x82_r_tb = 16'b1111111110100010;
   x82_i_tb = 16'b0;
   x83_r_tb = 16'b1111111110010000;
   x83_i_tb = 16'b0;
   x84_r_tb = 16'b1111111110010011;
   x84_i_tb = 16'b0;
   x85_r_tb = 16'b1111111110100001;
   x85_i_tb = 16'b0;
   x86_r_tb = 16'b1111111110101011;
   x86_i_tb = 16'b0;
   x87_r_tb = 16'b1111111110101100;
   x87_i_tb = 16'b0;
   x88_r_tb = 16'b1111111110101010;
   x88_i_tb = 16'b0;
   x89_r_tb = 16'b1111111110100111;
   x89_i_tb = 16'b0;
   x90_r_tb = 16'b1111111110101011;
   x90_i_tb = 16'b0;
   x91_r_tb = 16'b1111111110101100;
   x91_i_tb = 16'b0;
   x92_r_tb = 16'b1111111110101111;
   x92_i_tb = 16'b0;
   x93_r_tb = 16'b1111111110110000;
   x93_i_tb = 16'b0;
   x94_r_tb = 16'b1111111110101110;
   x94_i_tb = 16'b0;
   x95_r_tb = 16'b1111111110101010;
   x95_i_tb = 16'b0; 
    x96_r_tb = 16'b1111111110101000;
x96_i_tb =16'b0;
x97_r_tb = 16'b1111111110101100;
x97_i_tb =16'b0;
x98_r_tb = 16'b1111111110100111;
x98_i_tb =16'b0;
x99_r_tb = 16'b1111111110101010;
x99_i_tb =16'b0;
x100_r_tb = 16'b1111111110101011;
x100_i_tb =16'b0;
x101_r_tb = 16'b1111111110101010;
x101_i_tb =16'b0;
x102_r_tb = 16'b1111111110101011;
x102_i_tb =16'b0;
x103_r_tb = 16'b1111111110101100;
x103_i_tb =16'b0;
x104_r_tb = 16'b1111111110101011;
x104_i_tb =16'b0;
    x105_r_tb = 16'b1111111110101011;
   x105_i_tb = 16'b0;
   x106_r_tb = 16'b1111111110100111;
   x106_i_tb = 16'b0;
   x107_r_tb = 16'b1111111110100101;
   x107_i_tb = 16'b0;
   x108_r_tb = 16'b1111111110101010;
   x108_i_tb = 16'b0;
   x109_r_tb = 16'b1111111110101100;
   x109_i_tb = 16'b0;
   x110_r_tb = 16'b1111111110110001;
   x110_i_tb = 16'b0;
   x111_r_tb = 16'b1111111110101110;
   x111_i_tb = 16'b0;
   x112_r_tb = 16'b1111111110101110;
   x112_i_tb = 16'b0;
   x113_r_tb = 16'b1111111110101011;
   x113_i_tb = 16'b0;
   x114_r_tb = 16'b1111111110101000;
   x114_i_tb = 16'b0;
   x115_r_tb = 16'b1111111110101010;
   x115_i_tb = 16'b0;
   x116_r_tb = 16'b1111111110101000;
   x116_i_tb = 16'b0;
   x117_r_tb = 16'b1111111110100111;
   x117_i_tb = 16'b0;
   x118_r_tb = 16'b1111111110100101;
   x118_i_tb = 16'b0;
   x119_r_tb = 16'b1111111110100101;
   x119_i_tb = 16'b0;
   x120_r_tb = 16'b1111111110101000;
   x120_i_tb = 16'b0;
   x121_r_tb = 16'b1111111110101011;
   x121_i_tb = 16'b0;
   x122_r_tb = 16'b1111111110101011;
   x122_i_tb = 16'b0;
   x123_r_tb = 16'b1111111110101011;
   x123_i_tb = 16'b0;
   x124_r_tb = 16'b1111111110101000;
   x124_i_tb = 16'b0;
   x125_r_tb = 16'b1111111110100110;
   x125_i_tb = 16'b0;
   x126_r_tb = 16'b1111111110101100;
   x126_i_tb = 16'b0;
   x127_r_tb = 16'b1111111110101100;
   x127_i_tb = 16'b0; 
   ready_inputs_tb = 1'b1 ;
    #(4*Clock_Period)
   ready_inputs_tb = 1'b0 ;
   inputs = $fopen("inputs.txt", "r");

  end
endtask

task FFT_Operation;
begin
  wait(UUT_CWT_TOP.FFT.correct == 1) /* wait till the correct signal gets high then check the outputs */
  $display("X0 real is %b",UUT_CWT_TOP.FFT.X0_r);
end
endtask
endmodule