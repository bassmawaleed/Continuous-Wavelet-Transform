module IFFT_Time_Share_Top_Module_tb();
	
	
	/* Parameters */
	parameter Clock_Period = 4 ;
	parameter BITS =16;
	/* FIRST : Define the testbench signals */
	///////////// Inputs /////////////
    reg ready_inputs_tb ;
    reg clk_tb;
    reg rst_tb;
    reg [BITS-1 : 0 ] x0_r_tb ;
    reg [BITS-1 : 0 ] x0_i_tb ;
    reg [BITS-1 : 0 ] x1_r_tb ;
    reg [BITS-1 : 0 ] x1_i_tb ;
    reg [BITS-1 : 0 ] x2_r_tb ;
    reg [BITS-1 : 0 ] x2_i_tb;
    reg [BITS-1 : 0 ] x3_r_tb ;
    reg [BITS-1 : 0 ] x3_i_tb ;
    reg [BITS-1 : 0 ] x4_r_tb ;
    reg [BITS-1 : 0 ] x4_i_tb ;
    reg [BITS-1 : 0 ] x5_r_tb ;
    reg [BITS-1 : 0 ] x5_i_tb ;
    reg [BITS-1 : 0 ] x6_r_tb ;
    reg [BITS-1 : 0 ] x6_i_tb ;
    reg[BITS-1 : 0 ] x7_r_tb ;
    reg [BITS-1 : 0 ] x7_i_tb;
    reg [BITS-1 : 0 ] x8_r_tb;
    reg [BITS-1 : 0 ] x8_i_tb;
    reg [BITS-1 : 0 ] x9_r_tb;
    reg [BITS-1 : 0 ] x9_i_tb;
    reg [BITS-1 : 0 ] x10_r_tb;
    reg [BITS-1 : 0 ] x10_i_tb;
    reg [BITS-1 : 0 ] x11_r_tb;
    reg [BITS-1 : 0 ] x11_i_tb;
    reg [BITS-1 : 0 ] x12_r_tb;
    reg [BITS-1 : 0 ] x12_i_tb;
    reg [BITS-1 : 0 ] x13_r_tb;
    reg [BITS-1 : 0 ] x13_i_tb;
    reg [BITS-1 : 0 ] x14_r_tb;
    reg [BITS-1 : 0 ] x14_i_tb;
    reg [BITS-1 : 0 ] x15_r_tb;
    reg [BITS-1 : 0 ] x15_i_tb;
    reg [BITS-1 : 0 ] x16_r_tb ;
    reg [BITS-1 : 0 ] x16_i_tb ;
    reg [BITS-1 : 0 ] x17_r_tb ;
    reg [BITS-1 : 0 ] x17_i_tb ;
    reg [BITS-1 : 0 ] x18_r_tb ;
    reg [BITS-1 : 0 ] x18_i_tb;
    reg [BITS-1 : 0 ] x19_r_tb ;
    reg [BITS-1 : 0 ] x19_i_tb ;
    reg [BITS-1 : 0 ] x20_r_tb ;
    reg [BITS-1 : 0 ] x20_i_tb ;
    reg [BITS-1 : 0 ] x21_r_tb ;
    reg [BITS-1 : 0 ] x21_i_tb ;
    reg [BITS-1 : 0 ] x22_r_tb ;
    reg [BITS-1 : 0 ] x22_i_tb ;
    reg [BITS-1 : 0 ] x23_r_tb ;
    reg [BITS-1 : 0 ] x23_i_tb ;
    reg[BITS-1 : 0 ] x24_r_tb ;
    reg [BITS-1 : 0 ] x24_i_tb;
    reg [BITS-1 : 0 ] x25_r_tb;
    reg [BITS-1 : 0 ] x25_i_tb;
    reg [BITS-1 : 0 ] x26_r_tb;
    reg [BITS-1 : 0 ] x26_i_tb;
    reg [BITS-1 : 0 ] x27_r_tb;
    reg [BITS-1 : 0 ] x27_i_tb;
    reg [BITS-1 : 0 ] x28_r_tb;
    reg [BITS-1 : 0 ] x28_i_tb;
    reg [BITS-1 : 0 ] x29_r_tb;
    reg [BITS-1 : 0 ] x29_i_tb;
    reg [BITS-1 : 0 ] x30_r_tb;
    reg [BITS-1 : 0 ] x30_i_tb;
    reg [BITS-1 : 0 ] x31_r_tb;
    reg[BITS-1 : 0 ] x31_i_tb;
    reg [BITS-1 : 0 ] x32_r_tb;
    reg [BITS-1 : 0 ] x32_i_tb;
    reg [BITS-1 : 0 ] x33_r_tb ;
    reg [BITS-1 : 0 ] x33_i_tb ;
    reg [BITS-1 : 0 ] x34_r_tb ;
    reg [BITS-1 : 0 ] x34_i_tb ;
    reg [BITS-1 : 0 ] x35_r_tb ;
    reg [BITS-1 : 0 ] x35_i_tb;
    reg [BITS-1 : 0 ] x36_r_tb ;
    reg [BITS-1 : 0 ] x36_i_tb ;
    reg [BITS-1 : 0 ] x37_r_tb ;
    reg [BITS-1 : 0 ] x37_i_tb ;
    reg [BITS-1 : 0 ] x38_r_tb ;
    reg [BITS-1 : 0 ] x38_i_tb ;
    reg [BITS-1 : 0 ] x39_r_tb ;
    reg [BITS-1 : 0 ] x39_i_tb ;
    reg[BITS-1 : 0 ] x40_r_tb ;
    reg [BITS-1 : 0 ] x40_i_tb;
    reg [BITS-1 : 0 ] x41_r_tb;
    reg [BITS-1 : 0 ] x41_i_tb;
    reg [BITS-1 : 0 ] x42_r_tb;
    reg [BITS-1 : 0 ] x42_i_tb;
    reg [BITS-1 : 0 ] x43_r_tb;
    reg [BITS-1 : 0 ] x43_i_tb;
    reg [BITS-1 : 0 ] x44_r_tb;
    reg [BITS-1 : 0 ] x44_i_tb;
    reg [BITS-1 : 0 ] x45_r_tb;
    reg [BITS-1 : 0 ] x45_i_tb;
    reg [BITS-1 : 0 ] x46_r_tb;
    reg [BITS-1 : 0 ] x46_i_tb;
    reg [BITS-1 : 0 ] x47_r_tb;
    reg[BITS-1 : 0 ] x47_i_tb;
    reg [BITS-1 : 0 ] x48_r_tb;
    reg [BITS-1 : 0 ] x48_i_tb;
    reg [BITS-1 : 0 ] x49_r_tb ;
    reg [BITS-1 : 0 ] x49_i_tb ;
    reg [BITS-1 : 0 ] x50_r_tb ;
    reg [BITS-1 : 0 ] x50_i_tb ;
    reg [BITS-1 : 0 ] x51_r_tb ;
    reg [BITS-1 : 0 ] x51_i_tb;
    reg [BITS-1 : 0 ] x52_r_tb ;
    reg [BITS-1 : 0 ] x52_i_tb ;
    reg [BITS-1 : 0 ] x53_r_tb ;
    reg [BITS-1 : 0 ] x53_i_tb ;
    reg [BITS-1 : 0 ] x54_r_tb ;
    reg [BITS-1 : 0 ] x54_i_tb ;
    reg [BITS-1 : 0 ] x55_r_tb ;
    reg [BITS-1 : 0 ] x55_i_tb ;
    reg[BITS-1 : 0 ] x56_r_tb ;
    reg [BITS-1 : 0 ] x56_i_tb;
    reg [BITS-1 : 0 ] x57_r_tb;
    reg [BITS-1 : 0 ] x57_i_tb;
    reg [BITS-1 : 0 ] x58_r_tb;
    reg [BITS-1 : 0 ] x58_i_tb;
    reg [BITS-1 : 0 ] x59_r_tb;
    reg [BITS-1 : 0 ] x59_i_tb;
    reg [BITS-1 : 0 ] x60_r_tb;
    reg [BITS-1 : 0 ] x60_i_tb;
    reg [BITS-1 : 0 ] x61_r_tb;
    reg [BITS-1 : 0 ] x61_i_tb;
    reg [BITS-1 : 0 ] x62_r_tb;
    reg [BITS-1 : 0 ] x62_i_tb;
    reg [BITS-1 : 0 ] x63_r_tb;
    reg [BITS-1 : 0 ] x63_i_tb;
    reg [BITS-1 : 0 ] x64_r_tb;
    reg [BITS-1 : 0 ] x64_i_tb;
    reg [BITS-1 : 0 ] x65_r_tb ;
    reg [BITS-1 : 0 ] x65_i_tb ;
    reg [BITS-1 : 0 ] x66_r_tb ;
    reg [BITS-1 : 0 ] x66_i_tb ;
    reg [BITS-1 : 0 ] x67_r_tb ;
    reg [BITS-1 : 0 ] x67_i_tb;
    reg [BITS-1 : 0 ] x68_r_tb ;
    reg  [BITS-1 : 0 ] x68_i_tb ;
    reg [BITS-1 : 0 ] x69_r_tb ;
    reg [BITS-1 : 0 ] x69_i_tb ;
    reg [BITS-1 : 0 ] x70_r_tb ;
    reg [BITS-1 : 0 ] x70_i_tb ;
    reg [BITS-1 : 0 ] x71_r_tb ;
    reg [BITS-1 : 0 ] x71_i_tb ;
    reg [BITS-1 : 0 ] x72_r_tb ;
    reg [BITS-1 : 0 ] x72_i_tb;
    reg [BITS-1 : 0 ] x73_r_tb;
    reg [BITS-1 : 0 ] x73_i_tb;
    reg [BITS-1 : 0 ] x74_r_tb;
    reg [BITS-1 : 0 ] x74_i_tb;
    reg [BITS-1 : 0 ] x75_r_tb;
    reg [BITS-1 : 0 ] x75_i_tb;
    reg [BITS-1 : 0 ] x76_r_tb;
    reg [BITS-1 : 0 ] x76_i_tb;
    reg [BITS-1 : 0 ] x77_r_tb;
    reg [BITS-1 : 0 ] x77_i_tb;
    reg [BITS-1 : 0 ] x78_r_tb;
    reg [BITS-1 : 0 ] x78_i_tb;
    reg [BITS-1 : 0 ] x79_r_tb;
    reg [BITS-1 : 0 ] x79_i_tb;
    reg [BITS-1 : 0 ] x80_r_tb;
    reg [BITS-1 : 0 ] x80_i_tb;
    reg [BITS-1 : 0 ] x81_r_tb ;
    reg [BITS-1 : 0 ] x81_i_tb ;
    reg [BITS-1 : 0 ] x82_r_tb ;
    reg [BITS-1 : 0 ] x82_i_tb ;
    reg [BITS-1 : 0 ] x83_r_tb ;
    reg [BITS-1 : 0 ] x83_i_tb;
    reg [BITS-1 : 0 ] x84_r_tb ;
    reg [BITS-1 : 0 ] x84_i_tb ;
    reg [BITS-1 : 0 ] x85_r_tb ;
    reg [BITS-1 : 0 ] x85_i_tb ;
    reg [BITS-1 : 0 ] x86_r_tb ;
    reg [BITS-1 : 0 ] x86_i_tb ;
    reg [BITS-1 : 0 ] x87_r_tb ;
    reg [BITS-1 : 0 ] x87_i_tb ;
    reg[BITS-1 : 0 ] x88_r_tb ;
    reg [BITS-1 : 0 ] x88_i_tb;
    reg [BITS-1 : 0 ] x89_r_tb;
    reg [BITS-1 : 0 ] x89_i_tb;
    reg [BITS-1 : 0 ] x90_r_tb;
    reg [BITS-1 : 0 ] x90_i_tb;
    reg [BITS-1 : 0 ] x91_r_tb;
    reg [BITS-1 : 0 ] x91_i_tb;
    reg [BITS-1 : 0 ] x92_r_tb;
    reg [BITS-1 : 0 ] x92_i_tb;
    reg [BITS-1 : 0 ] x93_r_tb;
    reg [BITS-1 : 0 ] x93_i_tb;
    reg [BITS-1 : 0 ] x94_r_tb;
    reg [BITS-1 : 0 ] x94_i_tb;
    reg [BITS-1 : 0 ] x95_r_tb;
    reg [BITS-1 : 0 ] x95_i_tb;
    reg [BITS-1 : 0 ] x96_r_tb;
    reg [BITS-1 : 0 ] x96_i_tb;
    reg [BITS-1 : 0 ] x97_r_tb ;
    reg [BITS-1 : 0 ] x97_i_tb ;
    reg [BITS-1 : 0 ] x98_r_tb ;
    reg [BITS-1 : 0 ] x98_i_tb ;
    reg [BITS-1 : 0 ] x99_r_tb ;
    reg [BITS-1 : 0 ] x99_i_tb;
    reg [BITS-1 : 0 ] x100_r_tb ;
    reg [BITS-1 : 0 ] x100_i_tb ;
    reg [BITS-1 : 0 ] x101_r_tb ;
    reg [BITS-1 : 0 ] x101_i_tb ;
    reg [BITS-1 : 0 ] x102_r_tb ;
    reg [BITS-1 : 0 ] x102_i_tb ;
    reg [BITS-1 : 0 ] x103_r_tb ;
    reg [BITS-1 : 0 ] x103_i_tb ;
    reg [BITS-1 : 0 ] x104_r_tb ;
    reg [BITS-1 : 0 ] x104_i_tb;
    reg [BITS-1 : 0 ] x105_r_tb;
    reg [BITS-1 : 0 ] x105_i_tb;
    reg [BITS-1 : 0 ] x106_r_tb;
    reg [BITS-1 : 0 ] x106_i_tb;
    reg [BITS-1 : 0 ] x107_r_tb;
    reg [BITS-1 : 0 ] x107_i_tb;
    reg [BITS-1 : 0 ] x108_r_tb;
    reg [BITS-1 : 0 ] x108_i_tb;
    reg [BITS-1 : 0 ] x109_r_tb;
    reg [BITS-1 : 0 ] x109_i_tb;
    reg [BITS-1 : 0 ] x110_r_tb;
    reg [BITS-1 : 0 ] x110_i_tb;
    reg [BITS-1 : 0 ] x111_r_tb;
    reg [BITS-1 : 0 ] x111_i_tb;
    reg [BITS-1 : 0 ] x112_r_tb;
    reg [BITS-1 : 0 ] x112_i_tb;
    reg [BITS-1 : 0 ] x113_r_tb ;
    reg [BITS-1 : 0 ] x113_i_tb ;
    reg [BITS-1 : 0 ] x114_r_tb ;
    reg [BITS-1 : 0 ] x114_i_tb ;
    reg [BITS-1 : 0 ] x115_r_tb ;
    reg [BITS-1 : 0 ] x115_i_tb;
    reg [BITS-1 : 0 ] x116_r_tb ;
    reg [BITS-1 : 0 ] x116_i_tb ;
    reg [BITS-1 : 0 ] x117_r_tb ;
    reg [BITS-1 : 0 ] x117_i_tb ;
    reg [BITS-1 : 0 ] x118_r_tb ;
    reg [BITS-1 : 0 ] x118_i_tb ;
    reg [BITS-1 : 0 ] x119_r_tb ;
    reg [BITS-1 : 0 ] x119_i_tb ;
    reg [BITS-1 : 0 ] x120_r_tb ;
    reg [BITS-1 : 0 ] x120_i_tb;
    reg [BITS-1 : 0 ] x121_r_tb;
    reg [BITS-1 : 0 ] x121_i_tb;
    reg [BITS-1 : 0 ] x122_r_tb;
    reg [BITS-1 : 0 ] x122_i_tb;
    reg [BITS-1 : 0 ] x123_r_tb;
    reg [BITS-1 : 0 ] x123_i_tb;
    reg [BITS-1 : 0 ] x124_r_tb;
    reg [BITS-1 : 0 ] x124_i_tb;
    reg [BITS-1 : 0 ] x125_r_tb;
    reg [BITS-1 : 0 ] x125_i_tb;
    reg [BITS-1 : 0 ] x126_r_tb;
    reg [BITS-1 : 0 ] x126_i_tb;
    reg [BITS-1 : 0 ] x127_r_tb;
    reg [BITS-1 : 0 ] x127_i_tb;



    wire correct;
    wire [BITS-1 : 0 ] ifft_output0_r_tb;
    wire [BITS-1 : 0 ] ifft_output0_i_tb;
    wire [BITS-1 : 0 ] ifft_output1_r_tb;
    wire [BITS-1 : 0 ] ifft_output1_i_tb;
    wire [BITS-1 : 0 ] ifft_output2_r_tb;
    wire [BITS-1 : 0 ] ifft_output2_i_tb;
    wire [BITS-1 : 0 ] ifft_output3_r_tb;
    wire [BITS-1 : 0 ] ifft_output3_i_tb;
    wire [BITS-1 : 0 ] ifft_output4_r_tb;
    wire [BITS-1 : 0 ] ifft_output4_i_tb;
    wire [BITS-1 : 0 ] ifft_output5_r_tb;
    wire [BITS-1 : 0 ] ifft_output5_i_tb;
    wire [BITS-1 : 0 ] ifft_output6_r_tb;
    wire [BITS-1 : 0 ] ifft_output6_i_tb;
    wire [BITS-1 : 0 ] ifft_output7_r_tb;
    wire [BITS-1 : 0 ] ifft_output7_i_tb;
    wire [BITS-1 : 0 ] ifft_output8_r_tb;
    wire [BITS-1 : 0 ] ifft_output8_i_tb;
    wire [BITS-1 : 0 ] ifft_output9_r_tb;
    wire [BITS-1 : 0 ] ifft_output9_i_tb;
    wire [BITS-1 : 0 ] ifft_output10_r_tb;
    wire [BITS-1 : 0 ] ifft_output10_i_tb;
    wire [BITS-1 : 0 ] ifft_output11_r_tb;
    wire [BITS-1 : 0 ] ifft_output11_i_tb;
    wire [BITS-1 : 0 ] ifft_output12_r_tb;
    wire [BITS-1 : 0 ] ifft_output12_i_tb;
    wire [BITS-1 : 0 ] ifft_output13_r_tb;
    wire [BITS-1 : 0 ] ifft_output13_i_tb;
    wire [BITS-1 : 0 ] ifft_output14_r_tb;
    wire [BITS-1 : 0 ] ifft_output14_i_tb;
    wire [BITS-1 : 0 ] ifft_output15_r_tb;
    wire [BITS-1 : 0 ] ifft_output15_i_tb;
    wire [BITS-1 : 0 ] ifft_output16_r_tb;
    wire [BITS-1 : 0 ] ifft_output16_i_tb;
    wire [BITS-1 : 0 ] ifft_output17_r_tb;
    wire [BITS-1 : 0 ] ifft_output17_i_tb;
    wire [BITS-1 : 0 ] ifft_output18_r_tb;
    wire [BITS-1 : 0 ] ifft_output18_i_tb;
    wire [BITS-1 : 0 ] ifft_output19_r_tb;
    wire [BITS-1 : 0 ] ifft_output19_i_tb;
    wire [BITS-1 : 0 ] ifft_output20_r_tb;
    wire [BITS-1 : 0 ] ifft_output20_i_tb;
    wire [BITS-1 : 0 ] ifft_output21_r_tb;
    wire [BITS-1 : 0 ] ifft_output21_i_tb;
    wire [BITS-1 : 0 ] ifft_output22_r_tb;
    wire [BITS-1 : 0 ] ifft_output22_i_tb;
    wire [BITS-1 : 0 ] ifft_output23_r_tb;
    wire [BITS-1 : 0 ] ifft_output23_i_tb;
    wire [BITS-1 : 0 ] ifft_output24_r_tb;
    wire [BITS-1 : 0 ] ifft_output24_i_tb;
    wire [BITS-1 : 0 ] ifft_output25_r_tb;
    wire [BITS-1 : 0 ] ifft_output25_i_tb;
    wire [BITS-1 : 0 ] ifft_output26_r_tb;
    wire [BITS-1 : 0 ] ifft_output26_i_tb;
    wire [BITS-1 : 0 ] ifft_output27_r_tb;
    wire [BITS-1 : 0 ] ifft_output27_i_tb;
    wire [BITS-1 : 0 ] ifft_output28_r_tb;
    wire [BITS-1 : 0 ] ifft_output28_i_tb;
    wire [BITS-1 : 0 ] ifft_output29_r_tb;
    wire [BITS-1 : 0 ] ifft_output29_i_tb;
    wire [BITS-1 : 0 ] ifft_output30_r_tb;
    wire [BITS-1 : 0 ] ifft_output30_i_tb;
    wire [BITS-1 : 0 ] ifft_output31_r_tb;
    wire [BITS-1 : 0 ] ifft_output31_i_tb;
    wire [BITS-1 : 0 ] ifft_output32_r_tb;
    wire [BITS-1 : 0 ] ifft_output32_i_tb;
    wire [BITS-1 : 0 ] ifft_output33_r_tb;
    wire [BITS-1 : 0 ] ifft_output33_i_tb;
    wire [BITS-1 : 0 ] ifft_output34_r_tb;
    wire [BITS-1 : 0 ] ifft_output34_i_tb;
    wire [BITS-1 : 0 ] ifft_output35_r_tb;
    wire [BITS-1 : 0 ] ifft_output35_i_tb;
    wire [BITS-1 : 0 ] ifft_output36_r_tb;
    wire [BITS-1 : 0 ] ifft_output36_i_tb;
    wire [BITS-1 : 0 ] ifft_output37_r_tb;
    wire [BITS-1 : 0 ] ifft_output37_i_tb;
    wire [BITS-1 : 0 ] ifft_output38_r_tb;
    wire [BITS-1 : 0 ] ifft_output38_i_tb;
    wire [BITS-1 : 0 ] ifft_output39_r_tb;
    wire [BITS-1 : 0 ] ifft_output39_i_tb;
    wire [BITS-1 : 0 ] ifft_output40_r_tb;
    wire [BITS-1 : 0 ] ifft_output40_i_tb;
    wire [BITS-1 : 0 ] ifft_output41_r_tb;
    wire [BITS-1 : 0 ] ifft_output41_i_tb;
    wire [BITS-1 : 0 ] ifft_output42_r_tb;
    wire [BITS-1 : 0 ] ifft_output42_i_tb;
    wire [BITS-1 : 0 ] ifft_output43_r_tb;
    wire [BITS-1 : 0 ] ifft_output43_i_tb;
    wire [BITS-1 : 0 ] ifft_output44_r_tb;
    wire [BITS-1 : 0 ] ifft_output44_i_tb;
    wire [BITS-1 : 0 ] ifft_output45_r_tb;
    wire [BITS-1 : 0 ] ifft_output45_i_tb;
    wire [BITS-1 : 0 ] ifft_output46_r_tb;
    wire [BITS-1 : 0 ] ifft_output46_i_tb;
    wire [BITS-1 : 0 ] ifft_output47_r_tb;
    wire [BITS-1 : 0 ] ifft_output47_i_tb;
    wire [BITS-1 : 0 ] ifft_output48_r_tb;
    wire [BITS-1 : 0 ] ifft_output48_i_tb;
    wire [BITS-1 : 0 ] ifft_output49_r_tb;
    wire [BITS-1 : 0 ] ifft_output49_i_tb;
    wire [BITS-1 : 0 ] ifft_output50_r_tb;
    wire [BITS-1 : 0 ] ifft_output50_i_tb;
    wire [BITS-1 : 0 ] ifft_output51_r_tb;
    wire [BITS-1 : 0 ] ifft_output51_i_tb;
    wire [BITS-1 : 0 ] ifft_output52_r_tb;
    wire [BITS-1 : 0 ] ifft_output52_i_tb;
    wire [BITS-1 : 0 ] ifft_output53_r_tb;
    wire [BITS-1 : 0 ] ifft_output53_i_tb;
    wire [BITS-1 : 0 ] ifft_output54_r_tb;
    wire [BITS-1 : 0 ] ifft_output54_i_tb;
    wire [BITS-1 : 0 ] ifft_output55_r_tb;
    wire [BITS-1 : 0 ] ifft_output55_i_tb;
    wire [BITS-1 : 0 ] ifft_output56_r_tb;
    wire [BITS-1 : 0 ] ifft_output56_i_tb;
    wire [BITS-1 : 0 ] ifft_output57_r_tb;
    wire [BITS-1 : 0 ] ifft_output57_i_tb;
    wire [BITS-1 : 0 ] ifft_output58_r_tb;
    wire [BITS-1 : 0 ] ifft_output58_i_tb;
    wire [BITS-1 : 0 ] ifft_output59_r_tb;
    wire [BITS-1 : 0 ] ifft_output59_i_tb;
    wire [BITS-1 : 0 ] ifft_output60_r_tb;
    wire [BITS-1 : 0 ] ifft_output60_i_tb;
    wire [BITS-1 : 0 ] ifft_output61_r_tb;
    wire [BITS-1 : 0 ] ifft_output61_i_tb;
    wire [BITS-1 : 0 ] ifft_output62_r_tb;
    wire [BITS-1 : 0 ] ifft_output62_i_tb;
    wire [BITS-1 : 0 ] ifft_output63_r_tb;
    wire [BITS-1 : 0 ] ifft_output63_i_tb;
    wire [BITS-1 : 0 ] ifft_output64_r_tb;
    wire [BITS-1 : 0 ] ifft_output64_i_tb;
    wire [BITS-1 : 0 ] ifft_output65_r_tb;
    wire [BITS-1 : 0 ] ifft_output65_i_tb;
    wire [BITS-1 : 0 ] ifft_output66_r_tb;
    wire [BITS-1 : 0 ] ifft_output66_i_tb;
    wire [BITS-1 : 0 ] ifft_output67_r_tb;
    wire [BITS-1 : 0 ] ifft_output67_i_tb;
    wire [BITS-1 : 0 ] ifft_output68_r_tb;
    wire [BITS-1 : 0 ] ifft_output68_i_tb;
    wire [BITS-1 : 0 ] ifft_output69_r_tb;
    wire [BITS-1 : 0 ] ifft_output69_i_tb;
    wire [BITS-1 : 0 ] ifft_output70_r_tb;
    wire [BITS-1 : 0 ] ifft_output70_i_tb;
    wire [BITS-1 : 0 ] ifft_output71_r_tb;
    wire [BITS-1 : 0 ] ifft_output71_i_tb;
    wire [BITS-1 : 0 ] ifft_output72_r_tb;
    wire [BITS-1 : 0 ] ifft_output72_i_tb;
    wire [BITS-1 : 0 ] ifft_output73_r_tb;
    wire [BITS-1 : 0 ] ifft_output73_i_tb;
    wire [BITS-1 : 0 ] ifft_output74_r_tb;
    wire [BITS-1 : 0 ] ifft_output74_i_tb;
    wire [BITS-1 : 0 ] ifft_output75_r_tb;
    wire [BITS-1 : 0 ] ifft_output75_i_tb;
    wire [BITS-1 : 0 ] ifft_output76_r_tb;
    wire [BITS-1 : 0 ] ifft_output76_i_tb;
    wire [BITS-1 : 0 ] ifft_output77_r_tb;
    wire [BITS-1 : 0 ] ifft_output77_i_tb;
    wire [BITS-1 : 0 ] ifft_output78_r_tb;
    wire [BITS-1 : 0 ] ifft_output78_i_tb;
    wire [BITS-1 : 0 ] ifft_output79_r_tb;
    wire [BITS-1 : 0 ] ifft_output79_i_tb;
    wire [BITS-1 : 0 ] ifft_output80_r_tb;
    wire [BITS-1 : 0 ] ifft_output80_i_tb;
    wire [BITS-1 : 0 ] ifft_output81_r_tb;
    wire [BITS-1 : 0 ] ifft_output81_i_tb;
    wire [BITS-1 : 0 ] ifft_output82_r_tb;
    wire [BITS-1 : 0 ] ifft_output82_i_tb;
    wire [BITS-1 : 0 ] ifft_output83_r_tb;
    wire [BITS-1 : 0 ] ifft_output83_i_tb;
    wire [BITS-1 : 0 ] ifft_output84_r_tb;
    wire [BITS-1 : 0 ] ifft_output84_i_tb;
    wire [BITS-1 : 0 ] ifft_output85_r_tb;
    wire [BITS-1 : 0 ] ifft_output85_i_tb;
    wire [BITS-1 : 0 ] ifft_output86_r_tb;
    wire [BITS-1 : 0 ] ifft_output86_i_tb;
    wire [BITS-1 : 0 ] ifft_output87_r_tb;
    wire [BITS-1 : 0 ] ifft_output87_i_tb;
    wire [BITS-1 : 0 ] ifft_output88_r_tb;
    wire [BITS-1 : 0 ] ifft_output88_i_tb;
    wire [BITS-1 : 0 ] ifft_output89_r_tb;
    wire [BITS-1 : 0 ] ifft_output89_i_tb;
    wire [BITS-1 : 0 ] ifft_output90_r_tb;
    wire [BITS-1 : 0 ] ifft_output90_i_tb;
    wire [BITS-1 : 0 ] ifft_output91_r_tb;
    wire [BITS-1 : 0 ] ifft_output91_i_tb;
    wire [BITS-1 : 0 ] ifft_output92_r_tb;
    wire [BITS-1 : 0 ] ifft_output92_i_tb;
    wire [BITS-1 : 0 ] ifft_output93_r_tb;
    wire [BITS-1 : 0 ] ifft_output93_i_tb;
    wire [BITS-1 : 0 ] ifft_output94_r_tb;
    wire [BITS-1 : 0 ] ifft_output94_i_tb;
    wire [BITS-1 : 0 ] ifft_output95_r_tb;
    wire [BITS-1 : 0 ] ifft_output95_i_tb;
    wire [BITS-1 : 0 ] ifft_output96_r_tb;
    wire [BITS-1 : 0 ] ifft_output96_i_tb;
    wire [BITS-1 : 0 ] ifft_output97_r_tb;
    wire [BITS-1 : 0 ] ifft_output97_i_tb;
    wire [BITS-1 : 0 ] ifft_output98_r_tb;
    wire [BITS-1 : 0 ] ifft_output98_i_tb;
    wire [BITS-1 : 0 ] ifft_output99_r_tb;
    wire [BITS-1 : 0 ] ifft_output99_i_tb;
    wire [BITS-1 : 0 ] ifft_output100_r_tb;
    wire [BITS-1 : 0 ] ifft_output100_i_tb;
    wire [BITS-1 : 0 ] ifft_output101_r_tb;
    wire [BITS-1 : 0 ] ifft_output101_i_tb;
    wire [BITS-1 : 0 ] ifft_output102_r_tb;
    wire [BITS-1 : 0 ] ifft_output102_i_tb;
    wire [BITS-1 : 0 ] ifft_output103_r_tb;
    wire [BITS-1 : 0 ] ifft_output103_i_tb;
    wire [BITS-1 : 0 ] ifft_output104_r_tb;
    wire [BITS-1 : 0 ] ifft_output104_i_tb;
    wire [BITS-1 : 0 ] ifft_output105_r_tb;
    wire [BITS-1 : 0 ] ifft_output105_i_tb;
    wire [BITS-1 : 0 ] ifft_output106_r_tb;
    wire [BITS-1 : 0 ] ifft_output106_i_tb;
    wire [BITS-1 : 0 ] ifft_output107_r_tb;
    wire [BITS-1 : 0 ] ifft_output107_i_tb;
    wire [BITS-1 : 0 ] ifft_output108_r_tb;
    wire [BITS-1 : 0 ] ifft_output108_i_tb;
    wire [BITS-1 : 0 ] ifft_output109_r_tb;
    wire [BITS-1 : 0 ] ifft_output109_i_tb;
    wire [BITS-1 : 0 ] ifft_output110_r_tb;
    wire [BITS-1 : 0 ] ifft_output110_i_tb;
    wire [BITS-1 : 0 ] ifft_output111_r_tb;
    wire [BITS-1 : 0 ] ifft_output111_i_tb;
    wire [BITS-1 : 0 ] ifft_output112_r_tb;
    wire [BITS-1 : 0 ] ifft_output112_i_tb;
    wire [BITS-1 : 0 ] ifft_output113_r_tb;
    wire [BITS-1 : 0 ] ifft_output113_i_tb;
    wire [BITS-1 : 0 ] ifft_output114_r_tb;
    wire [BITS-1 : 0 ] ifft_output114_i_tb;
    wire [BITS-1 : 0 ] ifft_output115_r_tb;
    wire [BITS-1 : 0 ] ifft_output115_i_tb;
    wire [BITS-1 : 0 ] ifft_output116_r_tb;
    wire [BITS-1 : 0 ] ifft_output116_i_tb;
    wire [BITS-1 : 0 ] ifft_output117_r_tb;
    wire [BITS-1 : 0 ] ifft_output117_i_tb;
    wire [BITS-1 : 0 ] ifft_output118_r_tb;
    wire [BITS-1 : 0 ] ifft_output118_i_tb;
    wire [BITS-1 : 0 ] ifft_output119_r_tb;
    wire [BITS-1 : 0 ] ifft_output119_i_tb;
    wire [BITS-1 : 0 ] ifft_output120_r_tb;
    wire [BITS-1 : 0 ] ifft_output120_i_tb;
    wire [BITS-1 : 0 ] ifft_output121_r_tb;
    wire [BITS-1 : 0 ] ifft_output121_i_tb;
    wire [BITS-1 : 0 ] ifft_output122_r_tb;
    wire [BITS-1 : 0 ] ifft_output122_i_tb;
    wire [BITS-1 : 0 ] ifft_output123_r_tb;
    wire [BITS-1 : 0 ] ifft_output123_i_tb;
    wire [BITS-1 : 0 ] ifft_output124_r_tb;
    wire [BITS-1 : 0 ] ifft_output124_i_tb;
    wire [BITS-1 : 0 ] ifft_output125_r_tb;
    wire [BITS-1 : 0 ] ifft_output125_i_tb;
    wire [BITS-1 : 0 ] ifft_output126_r_tb;
    wire [BITS-1 : 0 ] ifft_output126_i_tb;
    wire [BITS-1 : 0 ] ifft_output127_r_tb;
    wire [BITS-1 : 0 ] ifft_output127_i_tb;


	/* SECOND : Instantiate the DesiXn Under Test */
	IFFT_Time_Share_Top_Module  DUT (
    .ready_inputs(ready_inputs_tb),
    .clk(clk_tb),
    .rst(rst_tb),
		.x0_r(x0_r_tb),
		.x0_i(x0_i_tb),
		.x1_r(x1_r_tb),
		.x1_i(x1_i_tb),
		.x2_r(x2_r_tb),
		.x2_i(x2_i_tb),
		.x3_r(x3_r_tb),
		.x3_i(x3_i_tb),
		.x4_r(x4_r_tb),
		.x4_i(x4_i_tb),
		.x5_r(x5_r_tb),
		.x5_i(x5_i_tb),
		.x6_r(x6_r_tb),
		.x6_i(x6_i_tb),
		.x7_r(x7_r_tb),
		.x7_i(x7_i_tb),
		.x8_r(x8_r_tb),
		.x8_i(x8_i_tb),
		.x9_r(x9_r_tb),
		.x9_i(x9_i_tb),
		.x10_r(x10_r_tb),
		.x10_i(x10_i_tb),
		.x11_r(x11_r_tb),
		.x11_i(x11_i_tb),
		.x12_r(x12_r_tb),
		.x12_i(x12_i_tb),
		.x13_r(x13_r_tb),
		.x13_i(x13_i_tb),
		.x14_r(x14_r_tb),
		.x14_i(x14_i_tb),
		.x15_r(x15_r_tb),
		.x15_i(x15_i_tb),
		.x16_r(x16_r_tb),
		.x16_i(x16_i_tb),
		.x17_r(x17_r_tb),
		.x17_i(x17_i_tb),
		.x18_r(x18_r_tb),
		.x18_i(x18_i_tb),
		.x19_r(x19_r_tb),
		.x19_i(x19_i_tb),
		.x20_r(x20_r_tb),
		.x20_i(x20_i_tb),
		.x21_r(x21_r_tb),
		.x21_i(x21_i_tb),
		.x22_r(x22_r_tb),
		.x22_i(x22_i_tb),
		.x23_r(x23_r_tb),
		.x23_i(x23_i_tb),
		.x24_r(x24_r_tb),
		.x24_i(x24_i_tb),
		.x25_r(x25_r_tb),
		.x25_i(x25_i_tb),
		.x26_r(x26_r_tb),
		.x26_i(x26_i_tb),
		.x27_r(x27_r_tb),
		.x27_i(x27_i_tb),
		.x28_r(x28_r_tb),
		.x28_i(x28_i_tb),
		.x29_r(x29_r_tb),
		.x29_i(x29_i_tb),
		.x30_r(x30_r_tb),
		.x30_i(x30_i_tb),
		.x31_r(x31_r_tb),
		.x31_i(x31_i_tb),
		.x32_r(x32_r_tb),
		.x32_i(x32_i_tb),
		.x33_r(x33_r_tb),
		.x33_i(x33_i_tb),
		.x34_r(x34_r_tb),
		.x34_i(x34_i_tb),
		.x35_r(x35_r_tb),
		.x35_i(x35_i_tb),
		.x36_r(x36_r_tb),
		.x36_i(x36_i_tb),
		.x37_r(x37_r_tb),
		.x37_i(x37_i_tb),
		.x38_r(x38_r_tb),
		.x38_i(x38_i_tb),
		.x39_r(x39_r_tb),
		.x39_i(x39_i_tb),
		.x40_r(x40_r_tb),
		.x40_i(x40_i_tb),
		.x41_r(x41_r_tb),
		.x41_i(x41_i_tb),
		.x42_r(x42_r_tb),
		.x42_i(x42_i_tb),
		.x43_r(x43_r_tb),
		.x43_i(x43_i_tb),
		.x44_r(x44_r_tb),
		.x44_i(x44_i_tb),
		.x45_r(x45_r_tb),
		.x45_i(x45_i_tb),
		.x46_r(x46_r_tb),
		.x46_i(x46_i_tb),
		.x47_r(x47_r_tb),
		.x47_i(x47_i_tb),
		.x48_r(x48_r_tb),
		.x48_i(x48_i_tb),
		.x49_r(x49_r_tb),
		.x49_i(x49_i_tb),
		.x50_r(x50_r_tb),
		.x50_i(x50_i_tb),
		.x51_r(x51_r_tb),
		.x51_i(x51_i_tb),
		.x52_r(x52_r_tb),
		.x52_i(x52_i_tb),
		.x53_r(x53_r_tb),
		.x53_i(x53_i_tb),
		.x54_r(x54_r_tb),
		.x54_i(x54_i_tb),
		.x55_r(x55_r_tb),
		.x55_i(x55_i_tb),
		.x56_r(x56_r_tb),
		.x56_i(x56_i_tb),
		.x57_r(x57_r_tb),
		.x57_i(x57_i_tb),
		.x58_r(x58_r_tb),
		.x58_i(x58_i_tb),
		.x59_r(x59_r_tb),
		.x59_i(x59_i_tb),
		.x60_r(x60_r_tb),
		.x60_i(x60_i_tb),
		.x61_r(x61_r_tb),
		.x61_i(x61_i_tb),
		.x62_r(x62_r_tb),
		.x62_i(x62_i_tb),
		.x63_r(x63_r_tb),
		.x63_i(x63_i_tb),
		.x64_r(x64_r_tb),
		.x64_i(x64_i_tb),
		.x65_r(x65_r_tb),
		.x65_i(x65_i_tb),
		.x66_r(x66_r_tb),
		.x66_i(x66_i_tb),
		.x67_r(x67_r_tb),
		.x67_i(x67_i_tb),
		.x68_r(x68_r_tb),
		.x68_i(x68_i_tb),
		.x69_r(x69_r_tb),
		.x69_i(x69_i_tb),
		.x70_r(x70_r_tb),
		.x70_i(x70_i_tb),
		.x71_r(x71_r_tb),
		.x71_i(x71_i_tb),
		.x72_r(x72_r_tb),
		.x72_i(x72_i_tb),
		.x73_r(x73_r_tb),
		.x73_i(x73_i_tb),
		.x74_r(x74_r_tb),
		.x74_i(x74_i_tb),
		.x75_r(x75_r_tb),
		.x75_i(x75_i_tb),
		.x76_r(x76_r_tb),
		.x76_i(x76_i_tb),
		.x77_r(x77_r_tb),
		.x77_i(x77_i_tb),
		.x78_r(x78_r_tb),
		.x78_i(x78_i_tb),
		.x79_r(x79_r_tb),
		.x79_i(x79_i_tb),
		.x80_r(x80_r_tb),
		.x80_i(x80_i_tb),
		.x81_r(x81_r_tb),
		.x81_i(x81_i_tb),
		.x82_r(x82_r_tb),
		.x82_i(x82_i_tb),
		.x83_r(x83_r_tb),
		.x83_i(x83_i_tb),
		.x84_r(x84_r_tb),
		.x84_i(x84_i_tb),
		.x85_r(x85_r_tb),
		.x85_i(x85_i_tb),
		.x86_r(x86_r_tb),
		.x86_i(x86_i_tb),
		.x87_r(x87_r_tb),
		.x87_i(x87_i_tb),
		.x88_r(x88_r_tb),
		.x88_i(x88_i_tb),
		.x89_r(x89_r_tb),
		.x89_i(x89_i_tb),
		.x90_r(x90_r_tb),
		.x90_i(x90_i_tb),
		.x91_r(x91_r_tb),
		.x91_i(x91_i_tb),
		.x92_r(x92_r_tb),
		.x92_i(x92_i_tb),
		.x93_r(x93_r_tb),
		.x93_i(x93_i_tb),
		.x94_r(x94_r_tb),
		.x94_i(x94_i_tb),
		.x95_r(x95_r_tb),
		.x95_i(x95_i_tb),
		.x96_r(x96_r_tb),
		.x96_i(x96_i_tb),
		.x97_r(x97_r_tb),
		.x97_i(x97_i_tb),
		.x98_r(x98_r_tb),
		.x98_i(x98_i_tb),
		.x99_r(x99_r_tb),
		.x99_i(x99_i_tb),
		.x100_r(x100_r_tb),
		.x100_i(x100_i_tb),
		.x101_r(x101_r_tb),
		.x101_i(x101_i_tb),
		.x102_r(x102_r_tb),
		.x102_i(x102_i_tb),
		.x103_r(x103_r_tb),
		.x103_i(x103_i_tb),
		.x104_r(x104_r_tb),
		.x104_i(x104_i_tb),
		.x105_r(x105_r_tb),
		.x105_i(x105_i_tb),
		.x106_r(x106_r_tb),
		.x106_i(x106_i_tb),
		.x107_r(x107_r_tb),
		.x107_i(x107_i_tb),
		.x108_r(x108_r_tb),
		.x108_i(x108_i_tb),
		.x109_r(x109_r_tb),
		.x109_i(x109_i_tb),
		.x110_r(x110_r_tb),
		.x110_i(x110_i_tb),
		.x111_r(x111_r_tb),
		.x111_i(x111_i_tb),
		.x112_r(x112_r_tb),
		.x112_i(x112_i_tb),
		.x113_r(x113_r_tb),
		.x113_i(x113_i_tb),
		.x114_r(x114_r_tb),
		.x114_i(x114_i_tb),
		.x115_r(x115_r_tb),
		.x115_i(x115_i_tb),
		.x116_r(x116_r_tb),
		.x116_i(x116_i_tb),
		.x117_r(x117_r_tb),
		.x117_i(x117_i_tb),
		.x118_r(x118_r_tb),
		.x118_i(x118_i_tb),
		.x119_r(x119_r_tb),
		.x119_i(x119_i_tb),
		.x120_r(x120_r_tb),
		.x120_i(x120_i_tb),
		.x121_r(x121_r_tb),
		.x121_i(x121_i_tb),
		.x122_r(x122_r_tb),
		.x122_i(x122_i_tb),
		.x123_r(x123_r_tb),
		.x123_i(x123_i_tb),
		.x124_r(x124_r_tb),
		.x124_i(x124_i_tb),
		.x125_r(x125_r_tb),
		.x125_i(x125_i_tb),
		.x126_r(x126_r_tb),
		.x126_i(x126_i_tb),
		.x127_r(x127_r_tb),
		.x127_i(x127_i_tb),
		


    .correct(correct),
    .ifft_output0_r(ifft_output0_r_tb),
    .ifft_output0_i(ifft_output0_i_tb),
    .ifft_output1_r(ifft_output1_r_tb),
    .ifft_output1_i(ifft_output1_i_tb),
    .ifft_output2_r(ifft_output2_r_tb),
    .ifft_output2_i(ifft_output2_i_tb),
    .ifft_output3_r(ifft_output3_r_tb),
    .ifft_output3_i(ifft_output3_i_tb),
    .ifft_output4_r(ifft_output4_r_tb),
    .ifft_output4_i(ifft_output4_i_tb),
    .ifft_output5_r(ifft_output5_r_tb),
    .ifft_output5_i(ifft_output5_i_tb),
    .ifft_output6_r(ifft_output6_r_tb),
    .ifft_output6_i(ifft_output6_i_tb),
    .ifft_output7_r(ifft_output7_r_tb),
    .ifft_output7_i(ifft_output7_i_tb),
    .ifft_output8_r(ifft_output8_r_tb),
    .ifft_output8_i(ifft_output8_i_tb),
    .ifft_output9_r(ifft_output9_r_tb),
    .ifft_output9_i(ifft_output9_i_tb),
    .ifft_output10_r(ifft_output10_r_tb),
    .ifft_output10_i(ifft_output10_i_tb),
    .ifft_output11_r(ifft_output11_r_tb),
    .ifft_output11_i(ifft_output11_i_tb),
    .ifft_output12_r(ifft_output12_r_tb),
    .ifft_output12_i(ifft_output12_i_tb),
    .ifft_output13_r(ifft_output13_r_tb),
    .ifft_output13_i(ifft_output13_i_tb),
    .ifft_output14_r(ifft_output14_r_tb),
    .ifft_output14_i(ifft_output14_i_tb),
    .ifft_output15_r(ifft_output15_r_tb),
    .ifft_output15_i(ifft_output15_i_tb),
    .ifft_output16_r(ifft_output16_r_tb),
    .ifft_output16_i(ifft_output16_i_tb),
    .ifft_output17_r(ifft_output17_r_tb),
    .ifft_output17_i(ifft_output17_i_tb),
    .ifft_output18_r(ifft_output18_r_tb),
    .ifft_output18_i(ifft_output18_i_tb),
    .ifft_output19_r(ifft_output19_r_tb),
    .ifft_output19_i(ifft_output19_i_tb),
    .ifft_output20_r(ifft_output20_r_tb),
    .ifft_output20_i(ifft_output20_i_tb),
    .ifft_output21_r(ifft_output21_r_tb),
    .ifft_output21_i(ifft_output21_i_tb),
    .ifft_output22_r(ifft_output22_r_tb),
    .ifft_output22_i(ifft_output22_i_tb),
    .ifft_output23_r(ifft_output23_r_tb),
    .ifft_output23_i(ifft_output23_i_tb),
    .ifft_output24_r(ifft_output24_r_tb),
    .ifft_output24_i(ifft_output24_i_tb),
    .ifft_output25_r(ifft_output25_r_tb),
    .ifft_output25_i(ifft_output25_i_tb),
    .ifft_output26_r(ifft_output26_r_tb),
    .ifft_output26_i(ifft_output26_i_tb),
    .ifft_output27_r(ifft_output27_r_tb),
    .ifft_output27_i(ifft_output27_i_tb),
    .ifft_output28_r(ifft_output28_r_tb),
    .ifft_output28_i(ifft_output28_i_tb),
    .ifft_output29_r(ifft_output29_r_tb),
    .ifft_output29_i(ifft_output29_i_tb),
    .ifft_output30_r(ifft_output30_r_tb),
    .ifft_output30_i(ifft_output30_i_tb),
    .ifft_output31_r(ifft_output31_r_tb),
    .ifft_output31_i(ifft_output31_i_tb),
    .ifft_output32_r(ifft_output32_r_tb),
    .ifft_output32_i(ifft_output32_i_tb),
    .ifft_output33_r(ifft_output33_r_tb),
    .ifft_output33_i(ifft_output33_i_tb),
    .ifft_output34_r(ifft_output34_r_tb),
    .ifft_output34_i(ifft_output34_i_tb),
    .ifft_output35_r(ifft_output35_r_tb),
    .ifft_output35_i(ifft_output35_i_tb),
    .ifft_output36_r(ifft_output36_r_tb),
    .ifft_output36_i(ifft_output36_i_tb),
    .ifft_output37_r(ifft_output37_r_tb),
    .ifft_output37_i(ifft_output37_i_tb),
    .ifft_output38_r(ifft_output38_r_tb),
    .ifft_output38_i(ifft_output38_i_tb),
    .ifft_output39_r(ifft_output39_r_tb),
    .ifft_output39_i(ifft_output39_i_tb),
    .ifft_output40_r(ifft_output40_r_tb),
    .ifft_output40_i(ifft_output40_i_tb),
    .ifft_output41_r(ifft_output41_r_tb),
    .ifft_output41_i(ifft_output41_i_tb),
    .ifft_output42_r(ifft_output42_r_tb),
    .ifft_output42_i(ifft_output42_i_tb),
    .ifft_output43_r(ifft_output43_r_tb),
    .ifft_output43_i(ifft_output43_i_tb),
    .ifft_output44_r(ifft_output44_r_tb),
    .ifft_output44_i(ifft_output44_i_tb),
    .ifft_output45_r(ifft_output45_r_tb),
    .ifft_output45_i(ifft_output45_i_tb),
    .ifft_output46_r(ifft_output46_r_tb),
    .ifft_output46_i(ifft_output46_i_tb),
    .ifft_output47_r(ifft_output47_r_tb),
    .ifft_output47_i(ifft_output47_i_tb),
    .ifft_output48_r(ifft_output48_r_tb),
    .ifft_output48_i(ifft_output48_i_tb),
    .ifft_output49_r(ifft_output49_r_tb),
    .ifft_output49_i(ifft_output49_i_tb),
    .ifft_output50_r(ifft_output50_r_tb),
    .ifft_output50_i(ifft_output50_i_tb),
    .ifft_output51_r(ifft_output51_r_tb),
    .ifft_output51_i(ifft_output51_i_tb),
    .ifft_output52_r(ifft_output52_r_tb),
    .ifft_output52_i(ifft_output52_i_tb),
    .ifft_output53_r(ifft_output53_r_tb),
    .ifft_output53_i(ifft_output53_i_tb),
    .ifft_output54_r(ifft_output54_r_tb),
    .ifft_output54_i(ifft_output54_i_tb),
    .ifft_output55_r(ifft_output55_r_tb),
    .ifft_output55_i(ifft_output55_i_tb),
    .ifft_output56_r(ifft_output56_r_tb),
    .ifft_output56_i(ifft_output56_i_tb),
    .ifft_output57_r(ifft_output57_r_tb),
    .ifft_output57_i(ifft_output57_i_tb),
    .ifft_output58_r(ifft_output58_r_tb),
    .ifft_output58_i(ifft_output58_i_tb),
    .ifft_output59_r(ifft_output59_r_tb),
    .ifft_output59_i(ifft_output59_i_tb),
    .ifft_output60_r(ifft_output60_r_tb),
    .ifft_output60_i(ifft_output60_i_tb),
    .ifft_output61_r(ifft_output61_r_tb),
    .ifft_output61_i(ifft_output61_i_tb),
    .ifft_output62_r(ifft_output62_r_tb),
    .ifft_output62_i(ifft_output62_i_tb),
    .ifft_output63_r(ifft_output63_r_tb),
    .ifft_output63_i(ifft_output63_i_tb),
    .ifft_output64_r(ifft_output64_r_tb),
    .ifft_output64_i(ifft_output64_i_tb),
    .ifft_output65_r(ifft_output65_r_tb),
    .ifft_output65_i(ifft_output65_i_tb),
    .ifft_output66_r(ifft_output66_r_tb),
    .ifft_output66_i(ifft_output66_i_tb),
    .ifft_output67_r(ifft_output67_r_tb),
    .ifft_output67_i(ifft_output67_i_tb),
    .ifft_output68_r(ifft_output68_r_tb),
    .ifft_output68_i(ifft_output68_i_tb),
    .ifft_output69_r(ifft_output69_r_tb),
    .ifft_output69_i(ifft_output69_i_tb),
    .ifft_output70_r(ifft_output70_r_tb),
    .ifft_output70_i(ifft_output70_i_tb),
    .ifft_output71_r(ifft_output71_r_tb),
    .ifft_output71_i(ifft_output71_i_tb),
    .ifft_output72_r(ifft_output72_r_tb),
    .ifft_output72_i(ifft_output72_i_tb),
    .ifft_output73_r(ifft_output73_r_tb),
    .ifft_output73_i(ifft_output73_i_tb),
    .ifft_output74_r(ifft_output74_r_tb),
    .ifft_output74_i(ifft_output74_i_tb),
    .ifft_output75_r(ifft_output75_r_tb),
    .ifft_output75_i(ifft_output75_i_tb),
    .ifft_output76_r(ifft_output76_r_tb),
    .ifft_output76_i(ifft_output76_i_tb),
    .ifft_output77_r(ifft_output77_r_tb),
    .ifft_output77_i(ifft_output77_i_tb),
    .ifft_output78_r(ifft_output78_r_tb),
    .ifft_output78_i(ifft_output78_i_tb),
    .ifft_output79_r(ifft_output79_r_tb),
    .ifft_output79_i(ifft_output79_i_tb),
    .ifft_output80_r(ifft_output80_r_tb),
    .ifft_output80_i(ifft_output80_i_tb),
    .ifft_output81_r(ifft_output81_r_tb),
    .ifft_output81_i(ifft_output81_i_tb),
    .ifft_output82_r(ifft_output82_r_tb),
    .ifft_output82_i(ifft_output82_i_tb),
    .ifft_output83_r(ifft_output83_r_tb),
    .ifft_output83_i(ifft_output83_i_tb),
    .ifft_output84_r(ifft_output84_r_tb),
    .ifft_output84_i(ifft_output84_i_tb),
    .ifft_output85_r(ifft_output85_r_tb),
    .ifft_output85_i(ifft_output85_i_tb),
    .ifft_output86_r(ifft_output86_r_tb),
    .ifft_output86_i(ifft_output86_i_tb),
    .ifft_output87_r(ifft_output87_r_tb),
    .ifft_output87_i(ifft_output87_i_tb),
    .ifft_output88_r(ifft_output88_r_tb),
    .ifft_output88_i(ifft_output88_i_tb),
    .ifft_output89_r(ifft_output89_r_tb),
    .ifft_output89_i(ifft_output89_i_tb),
    .ifft_output90_r(ifft_output90_r_tb),
    .ifft_output90_i(ifft_output90_i_tb),
    .ifft_output91_r(ifft_output91_r_tb),
    .ifft_output91_i(ifft_output91_i_tb),
    .ifft_output92_r(ifft_output92_r_tb),
    .ifft_output92_i(ifft_output92_i_tb),
    .ifft_output93_r(ifft_output93_r_tb),
    .ifft_output93_i(ifft_output93_i_tb),
    .ifft_output94_r(ifft_output94_r_tb),
    .ifft_output94_i(ifft_output94_i_tb),
    .ifft_output95_r(ifft_output95_r_tb),
    .ifft_output95_i(ifft_output95_i_tb),
    .ifft_output96_r(ifft_output96_r_tb),
    .ifft_output96_i(ifft_output96_i_tb),
    .ifft_output97_r(ifft_output97_r_tb),
    .ifft_output97_i(ifft_output97_i_tb),
    .ifft_output98_r(ifft_output98_r_tb),
    .ifft_output98_i(ifft_output98_i_tb),
    .ifft_output99_r(ifft_output99_r_tb),
    .ifft_output99_i(ifft_output99_i_tb),
    .ifft_output100_r(ifft_output100_r_tb),
    .ifft_output100_i(ifft_output100_i_tb),
    .ifft_output101_r(ifft_output101_r_tb),
    .ifft_output101_i(ifft_output101_i_tb),
    .ifft_output102_r(ifft_output102_r_tb),
    .ifft_output102_i(ifft_output102_i_tb),
    .ifft_output103_r(ifft_output103_r_tb),
    .ifft_output103_i(ifft_output103_i_tb),
    .ifft_output104_r(ifft_output104_r_tb),
    .ifft_output104_i(ifft_output104_i_tb),
    .ifft_output105_r(ifft_output105_r_tb),
    .ifft_output105_i(ifft_output105_i_tb),
    .ifft_output106_r(ifft_output106_r_tb),
    .ifft_output106_i(ifft_output106_i_tb),
    .ifft_output107_r(ifft_output107_r_tb),
    .ifft_output107_i(ifft_output107_i_tb),
    .ifft_output108_r(ifft_output108_r_tb),
    .ifft_output108_i(ifft_output108_i_tb),
    .ifft_output109_r(ifft_output109_r_tb),
    .ifft_output109_i(ifft_output109_i_tb),
    .ifft_output110_r(ifft_output110_r_tb),
    .ifft_output110_i(ifft_output110_i_tb),
    .ifft_output111_r(ifft_output111_r_tb),
    .ifft_output111_i(ifft_output111_i_tb),
    .ifft_output112_r(ifft_output112_r_tb),
    .ifft_output112_i(ifft_output112_i_tb),
    .ifft_output113_r(ifft_output113_r_tb),
    .ifft_output113_i(ifft_output113_i_tb),
    .ifft_output114_r(ifft_output114_r_tb),
    .ifft_output114_i(ifft_output114_i_tb),
    .ifft_output115_r(ifft_output115_r_tb),
    .ifft_output115_i(ifft_output115_i_tb),
    .ifft_output116_r(ifft_output116_r_tb),
    .ifft_output116_i(ifft_output116_i_tb),
    .ifft_output117_r(ifft_output117_r_tb),
    .ifft_output117_i(ifft_output117_i_tb),
    .ifft_output118_r(ifft_output118_r_tb),
    .ifft_output118_i(ifft_output118_i_tb),
    .ifft_output119_r(ifft_output119_r_tb),
    .ifft_output119_i(ifft_output119_i_tb),
    .ifft_output120_r(ifft_output120_r_tb),
    .ifft_output120_i(ifft_output120_i_tb),
    .ifft_output121_r(ifft_output121_r_tb),
    .ifft_output121_i(ifft_output121_i_tb),
    .ifft_output122_r(ifft_output122_r_tb),
    .ifft_output122_i(ifft_output122_i_tb),
    .ifft_output123_r(ifft_output123_r_tb),
    .ifft_output123_i(ifft_output123_i_tb),
    .ifft_output124_r(ifft_output124_r_tb),
    .ifft_output124_i(ifft_output124_i_tb),
    .ifft_output125_r(ifft_output125_r_tb),
    .ifft_output125_i(ifft_output125_i_tb),
    .ifft_output126_r(ifft_output126_r_tb),
    .ifft_output126_i(ifft_output126_i_tb),
    .ifft_output127_r(ifft_output127_r_tb),
    .ifft_output127_i(ifft_output127_i_tb)
	);
	
	/* THIRD : Clock SiXnal Xeneration */
	always #(Clock_Period / 2) clk_tb = ~clk_tb ;
	
	/* FOURTH : Initial Block */
	initial begin
	$dumpfile("FFT_Time_Share.vcd");
	$dumpvars;

	initialize();

 
	reset();
  
	/* TEST CASE 1 */
	//TEST_CASE_1();
	
	TEST_CASE_1();
	

	
	
	#(100 * Clock_Period)
	$stop ;

end

task initialize ;
begin
  ready_inputs_tb = 1'b0;
  clk_tb = 1'b1 ; 
  rst_tb = 0;
x0_r_tb = 16'b00000000_00000000;
x0_i_tb = 16'b00000000_00000000;
x1_r_tb = 16'b00000000_00000000;
x1_i_tb = 16'b00000000_00000000;
x2_r_tb = 16'b00000000_00000000;
x2_i_tb = 16'b00000000_00000000;
x3_r_tb = 16'b00000000_00000000;
x3_i_tb = 16'b00000000_00000000;
x4_r_tb = 16'b00000000_00000000;
x4_i_tb = 16'b00000000_00000000;
x5_r_tb = 16'b00000000_00000000;
x5_i_tb = 16'b00000000_00000000;
x6_r_tb = 16'b00000000_00000000;
x6_i_tb = 16'b00000000_00000000;
x7_r_tb = 16'b00000000_00000000;
x7_i_tb = 16'b00000000_00000000;
x8_r_tb = 16'b00000000_00000000;
x8_i_tb = 16'b00000000_00000000;
x9_r_tb = 16'b00000000_00000000;
x9_i_tb = 16'b00000000_00000000;
x10_r_tb = 16'b00000000_00000000;
x10_i_tb = 16'b00000000_00000000;
x11_r_tb = 16'b00000000_00000000;
x11_i_tb = 16'b00000000_00000000;
x12_r_tb = 16'b00000000_00000000;
x12_i_tb = 16'b00000000_00000000;
x13_r_tb = 16'b00000000_00000000;
x13_i_tb = 16'b00000000_00000000;
x14_r_tb = 16'b00000000_00000000;
x14_i_tb = 16'b00000000_00000000;
x15_r_tb = 16'b00000000_00000000;
x15_i_tb = 16'b00000000_00000000;
x16_r_tb = 16'b00000000_00000000;
x16_i_tb = 16'b00000000_00000000;
x17_r_tb = 16'b00000000_00000000;
x17_i_tb = 16'b00000000_00000000;
x18_r_tb = 16'b00000000_00000000;
x18_i_tb = 16'b00000000_00000000;
x19_r_tb = 16'b00000000_00000000;
x19_i_tb = 16'b00000000_00000000;
x20_r_tb = 16'b00000000_00000000;
x20_i_tb = 16'b00000000_00000000;
x21_r_tb = 16'b00000000_00000000;
x21_i_tb = 16'b00000000_00000000;
x22_r_tb = 16'b00000000_00000000;
x22_i_tb = 16'b00000000_00000000;
x23_r_tb = 16'b00000000_00000000;
x23_i_tb = 16'b00000000_00000000;
x24_r_tb = 16'b00000000_00000000;
x24_i_tb = 16'b00000000_00000000;
x25_r_tb = 16'b00000000_00000000;
x25_i_tb = 16'b00000000_00000000;
x26_r_tb = 16'b00000000_00000000;
x26_i_tb = 16'b00000000_00000000;
x27_r_tb = 16'b00000000_00000000;
x27_i_tb = 16'b00000000_00000000;
x28_r_tb = 16'b00000000_00000000;
x28_i_tb = 16'b00000000_00000000;
x29_r_tb = 16'b00000000_00000000;
x29_i_tb = 16'b00000000_00000000;
x30_r_tb = 16'b00000000_00000000;
x30_i_tb = 16'b00000000_00000000;
x31_r_tb = 16'b00000000_00000000;
x31_i_tb = 16'b00000000_00000000;
x32_r_tb = 16'b00000000_00000000;
x32_i_tb = 16'b00000000_00000000;
x33_r_tb = 16'b00000000_00000000;
x33_i_tb = 16'b00000000_00000000;
x34_r_tb = 16'b00000000_00000000;
x34_i_tb = 16'b00000000_00000000;
x35_r_tb = 16'b00000000_00000000;
x35_i_tb = 16'b00000000_00000000;
x36_r_tb = 16'b00000000_00000000;
x36_i_tb = 16'b00000000_00000000;
x37_r_tb = 16'b00000000_00000000;
x37_i_tb = 16'b00000000_00000000;
x38_r_tb = 16'b00000000_00000000;
x38_i_tb = 16'b00000000_00000000;
x39_r_tb = 16'b00000000_00000000;
x39_i_tb = 16'b00000000_00000000;
x40_r_tb = 16'b00000000_00000000;
x40_i_tb = 16'b00000000_00000000;
x41_r_tb = 16'b00000000_00000000;
x41_i_tb = 16'b00000000_00000000;
x42_r_tb = 16'b00000000_00000000;
x42_i_tb = 16'b00000000_00000000;
x43_r_tb = 16'b00000000_00000000;
x43_i_tb = 16'b00000000_00000000;
x44_r_tb = 16'b00000000_00000000;
x44_i_tb = 16'b00000000_00000000;
x45_r_tb = 16'b00000000_00000000;
x45_i_tb = 16'b00000000_00000000;
x46_r_tb = 16'b00000000_00000000;
x46_i_tb = 16'b00000000_00000000;
x47_r_tb = 16'b00000000_00000000;
x47_i_tb = 16'b00000000_00000000;
x48_r_tb = 16'b00000000_00000000;
x48_i_tb = 16'b00000000_00000000;
x49_r_tb = 16'b00000000_00000000;
x49_i_tb = 16'b00000000_00000000;
x50_r_tb = 16'b00000000_00000000;
x50_i_tb = 16'b00000000_00000000;
x51_r_tb = 16'b00000000_00000000;
x51_i_tb = 16'b00000000_00000000;
x52_r_tb = 16'b00000000_00000000;
x52_i_tb = 16'b00000000_00000000;
x53_r_tb = 16'b00000000_00000000;
x53_i_tb = 16'b00000000_00000000;
x54_r_tb = 16'b00000000_00000000;
x54_i_tb = 16'b00000000_00000000;
x55_r_tb = 16'b00000000_00000000;
x55_i_tb = 16'b00000000_00000000;
x56_r_tb = 16'b00000000_00000000;
x56_i_tb = 16'b00000000_00000000;
x57_r_tb = 16'b00000000_00000000;
x57_i_tb = 16'b00000000_00000000;
x58_r_tb = 16'b00000000_00000000;
x58_i_tb = 16'b00000000_00000000;
x59_r_tb = 16'b00000000_00000000;
x59_i_tb = 16'b00000000_00000000;
x60_r_tb = 16'b00000000_00000000;
x60_i_tb = 16'b00000000_00000000;
x61_r_tb = 16'b00000000_00000000;
x61_i_tb = 16'b00000000_00000000;
x62_r_tb = 16'b00000000_00000000;
x62_i_tb = 16'b00000000_00000000;
x63_r_tb = 16'b00000000_00000000;
x63_i_tb = 16'b00000000_00000000;
x64_r_tb = 16'b00000000_00000000;
x64_i_tb = 16'b00000000_00000000;
x65_r_tb = 16'b00000000_00000000;
x65_i_tb = 16'b00000000_00000000;
x66_r_tb = 16'b00000000_00000000;
x66_i_tb = 16'b00000000_00000000;
x67_r_tb = 16'b00000000_00000000;
x67_i_tb = 16'b00000000_00000000;
x68_r_tb = 16'b00000000_00000000;
x68_i_tb = 16'b00000000_00000000;
x69_r_tb = 16'b00000000_00000000;
x69_i_tb = 16'b00000000_00000000;
x70_r_tb = 16'b00000000_00000000;
x70_i_tb = 16'b00000000_00000000;
x71_r_tb = 16'b00000000_00000000;
x71_i_tb = 16'b00000000_00000000;
x72_r_tb = 16'b00000000_00000000;
x72_i_tb = 16'b00000000_00000000;
x73_r_tb = 16'b00000000_00000000;
x73_i_tb = 16'b00000000_00000000;
x74_r_tb = 16'b00000000_00000000;
x74_i_tb = 16'b00000000_00000000;
x75_r_tb = 16'b00000000_00000000;
x75_i_tb = 16'b00000000_00000000;
x76_r_tb = 16'b00000000_00000000;
x76_i_tb = 16'b00000000_00000000;
x77_r_tb = 16'b00000000_00000000;
x77_i_tb = 16'b00000000_00000000;
x78_r_tb = 16'b00000000_00000000;
x78_i_tb = 16'b00000000_00000000;
x79_r_tb = 16'b00000000_00000000;
x79_i_tb = 16'b00000000_00000000;
x80_r_tb = 16'b00000000_00000000;
x80_i_tb = 16'b00000000_00000000;
x81_r_tb = 16'b00000000_00000000;
x81_i_tb = 16'b00000000_00000000;
x82_r_tb = 16'b00000000_00000000;
x82_i_tb = 16'b00000000_00000000;
x83_r_tb = 16'b00000000_00000000;
x83_i_tb = 16'b00000000_00000000;
x84_r_tb = 16'b00000000_00000000;
x84_i_tb = 16'b00000000_00000000;
x85_r_tb = 16'b00000000_00000000;
x85_i_tb = 16'b00000000_00000000;
x86_r_tb = 16'b00000000_00000000;
x86_i_tb = 16'b00000000_00000000;
x87_r_tb = 16'b00000000_00000000;
x87_i_tb = 16'b00000000_00000000;
x88_r_tb = 16'b00000000_00000000;
x88_i_tb = 16'b00000000_00000000;
x89_r_tb = 16'b00000000_00000000;
x89_i_tb = 16'b00000000_00000000;
x90_r_tb = 16'b00000000_00000000;
x90_i_tb = 16'b00000000_00000000;
x91_r_tb = 16'b00000000_00000000;
x91_i_tb = 16'b00000000_00000000;
x92_r_tb = 16'b00000000_00000000;
x92_i_tb = 16'b00000000_00000000;
x93_r_tb = 16'b00000000_00000000;
x93_i_tb = 16'b00000000_00000000;
x94_r_tb = 16'b00000000_00000000;
x94_i_tb = 16'b00000000_00000000;
x95_r_tb = 16'b00000000_00000000;
x95_i_tb = 16'b00000000_00000000;
x96_r_tb = 16'b00000000_00000000;
x96_i_tb = 16'b00000000_00000000;
x97_r_tb = 16'b00000000_00000000;
x97_i_tb = 16'b00000000_00000000;
x98_r_tb = 16'b00000000_00000000;
x98_i_tb = 16'b00000000_00000000;
x99_r_tb = 16'b00000000_00000000;
x99_i_tb = 16'b00000000_00000000;
x100_r_tb = 16'b00000000_00000000;
x100_i_tb = 16'b00000000_00000000;
x101_r_tb = 16'b00000000_00000000;
x101_i_tb = 16'b00000000_00000000;
x102_r_tb = 16'b00000000_00000000;
x102_i_tb = 16'b00000000_00000000;
x103_r_tb = 16'b00000000_00000000;
x103_i_tb = 16'b00000000_00000000;
x104_r_tb = 16'b00000000_00000000;
x104_i_tb = 16'b00000000_00000000;
x105_r_tb = 16'b00000000_00000000;
x105_i_tb = 16'b00000000_00000000;
x106_r_tb = 16'b00000000_00000000;
x106_i_tb = 16'b00000000_00000000;
x107_r_tb = 16'b00000000_00000000;
x107_i_tb = 16'b00000000_00000000;
x108_r_tb = 16'b00000000_00000000;
x108_i_tb = 16'b00000000_00000000;
x109_r_tb = 16'b00000000_00000000;
x109_i_tb = 16'b00000000_00000000;
x110_r_tb = 16'b00000000_00000000;
x110_i_tb = 16'b00000000_00000000;
x111_r_tb = 16'b00000000_00000000;
x111_i_tb = 16'b00000000_00000000;
x112_r_tb = 16'b00000000_00000000;
x112_i_tb = 16'b00000000_00000000;
x113_r_tb = 16'b00000000_00000000;
x113_i_tb = 16'b00000000_00000000;
x114_r_tb = 16'b00000000_00000000;
x114_i_tb = 16'b00000000_00000000;
x115_r_tb = 16'b00000000_00000000;
x115_i_tb = 16'b00000000_00000000;
x116_r_tb = 16'b00000000_00000000;
x116_i_tb = 16'b00000000_00000000;
x117_r_tb = 16'b00000000_00000000;
x117_i_tb = 16'b00000000_00000000;
x118_r_tb = 16'b00000000_00000000;
x118_i_tb = 16'b00000000_00000000;
x119_r_tb = 16'b00000000_00000000;
x119_i_tb = 16'b00000000_00000000;
x120_r_tb = 16'b00000000_00000000;
x120_i_tb = 16'b00000000_00000000;
x121_r_tb = 16'b00000000_00000000;
x121_i_tb = 16'b00000000_00000000;
x122_r_tb = 16'b00000000_00000000;
x122_i_tb = 16'b00000000_00000000;
x123_r_tb = 16'b00000000_00000000;
x123_i_tb = 16'b00000000_00000000;
x124_r_tb = 16'b00000000_00000000;
x124_i_tb = 16'b00000000_00000000;
x125_r_tb = 16'b00000000_00000000;
x125_i_tb = 16'b00000000_00000000;
x126_r_tb = 16'b00000000_00000000;
x126_i_tb = 16'b00000000_00000000;
x127_r_tb = 16'b00000000_00000000;
x127_i_tb = 16'b00000000_00000000;
end
endtask

task reset ;
  begin
	/* Reset */
    #(Clock_Period)
    rst_tb = 1'b1 ;
  end
endtask



task TEST_CASE_1;
  begin
	/* TEST CASE 2 */
  x0_r_tb = 16'b11111111_11011011;
x0_i_tb =16'b11111111_11110000;
x1_r_tb = 16'b11111111_11011011;
x1_i_tb =16'b11111111_11110000;
x2_r_tb = 16'b11111111_11011011;
x2_i_tb =16'b11111111_11110000;
x3_r_tb = 16'b11111111_11011011;
x3_i_tb =16'b11111111_11110000;
x4_r_tb = 16'b11111111_11011011;
x4_i_tb =16'b11111111_11110000;
x5_r_tb = 16'b11111111_11011011;
x5_i_tb =16'b11111111_11110000;
x6_r_tb = 16'b11111111_11011011;
x6_i_tb =16'b11111111_11110000;
x7_r_tb = 16'b11111111_11011011;
x7_i_tb =16'b11111111_11110000;
x8_r_tb = 16'b11111111_11011011;
x8_i_tb =16'b11111111_11110000;
    x9_r_tb = 16'b11111111_11100010;
   x9_i_tb = 16'b00000000_00010100;
   x10_r_tb = 16'b00000000_00100010;
   x10_i_tb = 16'b00000000_00010100;
   x11_r_tb = 16'b11111111_11011011;
   x11_i_tb = 16'b11111111_11101011;
   x12_r_tb = 16'b00000000_00100110;
   x12_i_tb = 16'b11111111_11101011;
   x13_r_tb = 16'b11111111_11011000;
   x13_i_tb = 16'b00000000_00010011;
   x14_r_tb = 16'b00000000_00100111;
   x14_i_tb = 16'b00000000_00010001;
   x15_r_tb = 16'b00000000_00101000;
   x15_i_tb = 16'b00000000_00010001;
   x16_r_tb = 16'b11111111_11010100;
   x16_i_tb = 16'b11111111_11110000;
   x17_r_tb = 16'b00000000_00101110;
   x17_i_tb = 16'b11111111_11110010;
   x18_r_tb = 16'b11111111_11010001;
   x18_i_tb = 16'b00000000_00001100;
   x19_r_tb = 16'b00000000_00101011;
   x19_i_tb = 16'b00000000_00001100;
   x20_r_tb = 16'b00000000_00100111;
   x20_i_tb = 16'b00000000_00001010;
   x21_r_tb = 16'b11111111_11010100;
   x21_i_tb = 16'b00000000_00001010;
   x22_r_tb = 16'b11111111_11010010;
   x22_i_tb = 16'b11111111_11110010;
   x23_r_tb = 16'b00000000_00110000;
   x23_i_tb = 16'b11111111_11101101;
   x24_r_tb = 16'b11111111_11010010;
   x24_i_tb = 16'b00000000_00010100;
   x25_r_tb = 16'b00000000_00100111;
   x25_i_tb = 16'b11111111_11101011;
   x26_r_tb = 16'b00000000_00100010;
   x26_i_tb = 16'b00000000_00010001;
   x27_r_tb = 16'b00000000_00100111;
   x27_i_tb = 16'b00000000_00010100;
   x28_r_tb = 16'b00000000_00110000;
   x28_i_tb = 16'b11111111_11101100;
   x29_r_tb = 16'b11111111_11001100;
   x29_i_tb = 16'b00000000_00010111;
   x30_r_tb = 16'b00000000_00111100;
   x30_i_tb = 16'b00000000_00011000;
   x31_r_tb = 16'b11111111_11000111;
   x31_i_tb = 16'b00000000_00010111; 
    x32_r_tb = 16'b11111111_11011011;
x32_i_tb =16'b11111111_11110000;
x33_r_tb = 16'b11111111_11011011;
x33_i_tb =16'b11111111_11110000;
x34_r_tb = 16'b11111111_11011011;
x34_i_tb =16'b11111111_11110000;
x35_r_tb = 16'b11111111_11011011;
x35_i_tb =16'b11111111_11110000;
x36_r_tb = 16'b11111111_11011011;
x36_i_tb =16'b11111111_11110000;
x37_r_tb = 16'b11111111_11011011;
x37_i_tb =16'b11111111_11110000;
x38_r_tb = 16'b11111111_11011011;
x38_i_tb =16'b11111111_11110000;
x39_r_tb = 16'b11111111_11011011;
x39_i_tb =16'b11111111_11110000;
x40_r_tb = 16'b11111111_11011011;
x40_i_tb =16'b11111111_11110000;
    x41_r_tb = 16'b11111111_11100010;
   x41_i_tb = 16'b00000000_00010100;
   x42_r_tb = 16'b00000000_00100010;
   x42_i_tb = 16'b00000000_00010100;
   x43_r_tb = 16'b11111111_11011011;
   x43_i_tb = 16'b11111111_11101011;
   x44_r_tb = 16'b00000000_00100110;
   x44_i_tb = 16'b11111111_11101011;
   x45_r_tb = 16'b11111111_11011000;
   x45_i_tb = 16'b00000000_00010011;
   x46_r_tb = 16'b00000000_00100111;
   x46_i_tb = 16'b00000000_00010001;
   x47_r_tb = 16'b00000000_00101000;
   x47_i_tb = 16'b00000000_00010001;
   x48_r_tb = 16'b11111111_11010100;
   x48_i_tb = 16'b11111111_11110000;
   x49_r_tb = 16'b00000000_00101110;
   x49_i_tb = 16'b11111111_11110010;
   x50_r_tb = 16'b11111111_11010001;
   x50_i_tb = 16'b00000000_00001100;
   x51_r_tb = 16'b00000000_00101011;
   x51_i_tb = 16'b00000000_00001100;
   x52_r_tb = 16'b00000000_00100111;
   x52_i_tb = 16'b00000000_00001010;
   x53_r_tb = 16'b11111111_11010100;
   x53_i_tb = 16'b00000000_00001010;
   x54_r_tb = 16'b11111111_11010010;
   x54_i_tb = 16'b11111111_11110010;
   x55_r_tb = 16'b00000000_00110000;
   x55_i_tb = 16'b11111111_11101101;
   x56_r_tb = 16'b11111111_11010010;
   x56_i_tb = 16'b00000000_00010100;
   x57_r_tb = 16'b00000000_00100111;
   x57_i_tb = 16'b11111111_11101011;
   x58_r_tb = 16'b00000000_00100010;
   x58_i_tb = 16'b00000000_00010001;
   x59_r_tb = 16'b00000000_00100111;
   x59_i_tb = 16'b00000000_00010100;
   x60_r_tb = 16'b00000000_00110000;
   x60_i_tb = 16'b11111111_11101100;
   x61_r_tb = 16'b11111111_11001100;
   x61_i_tb = 16'b00000000_00010111;
   x62_r_tb = 16'b00000000_00111100;
   x62_i_tb = 16'b00000000_00011000;
   x63_r_tb = 16'b11111111_11000111;
   x63_i_tb = 16'b00000000_00010111; 
    x64_r_tb = 16'b11111111_11011011;
x64_i_tb =16'b11111111_11110000;
x65_r_tb = 16'b11111111_11011011;
x65_i_tb =16'b11111111_11110000;
x66_r_tb = 16'b11111111_11011011;
x66_i_tb =16'b11111111_11110000;
x67_r_tb = 16'b11111111_11011011;
x67_i_tb =16'b11111111_11110000;
x68_r_tb = 16'b11111111_11011011;
x68_i_tb =16'b11111111_11110000;
x69_r_tb = 16'b11111111_11011011;
x69_i_tb =16'b11111111_11110000;
x70_r_tb = 16'b11111111_11011011;
x70_i_tb =16'b11111111_11110000;
x71_r_tb = 16'b11111111_11011011;
x71_i_tb =16'b11111111_11110000;
x72_r_tb = 16'b11111111_11011011;
x72_i_tb =16'b11111111_11110000;
    x73_r_tb = 16'b11111111_11100010;
   x73_i_tb = 16'b00000000_00010100;
   x74_r_tb = 16'b00000000_00100010;
   x74_i_tb = 16'b00000000_00010100;
   x75_r_tb = 16'b11111111_11011011;
   x75_i_tb = 16'b11111111_11101011;
   x76_r_tb = 16'b00000000_00100110;
   x76_i_tb = 16'b11111111_11101011;
   x77_r_tb = 16'b11111111_11011000;
   x77_i_tb = 16'b00000000_00010011;
   x78_r_tb = 16'b00000000_00100111;
   x78_i_tb = 16'b00000000_00010001;
   x79_r_tb = 16'b00000000_00101000;
   x79_i_tb = 16'b00000000_00010001;
   x80_r_tb = 16'b11111111_11010100;
   x80_i_tb = 16'b11111111_11110000;
   x81_r_tb = 16'b00000000_00101110;
   x81_i_tb = 16'b11111111_11110010;
   x82_r_tb = 16'b11111111_11010001;
   x82_i_tb = 16'b00000000_00001100;
   x83_r_tb = 16'b00000000_00101011;
   x83_i_tb = 16'b00000000_00001100;
   x84_r_tb = 16'b00000000_00100111;
   x84_i_tb = 16'b00000000_00001010;
   x85_r_tb = 16'b11111111_11010100;
   x85_i_tb = 16'b00000000_00001010;
   x86_r_tb = 16'b11111111_11010010;
   x86_i_tb = 16'b11111111_11110010;
   x87_r_tb = 16'b00000000_00110000;
   x87_i_tb = 16'b11111111_11101101;
   x88_r_tb = 16'b11111111_11010010;
   x88_i_tb = 16'b00000000_00010100;
   x89_r_tb = 16'b00000000_00100111;
   x89_i_tb = 16'b11111111_11101011;
   x90_r_tb = 16'b00000000_00100010;
   x90_i_tb = 16'b00000000_00010001;
   x91_r_tb = 16'b00000000_00100111;
   x91_i_tb = 16'b00000000_00010100;
   x92_r_tb = 16'b00000000_00110000;
   x92_i_tb = 16'b11111111_11101100;
   x93_r_tb = 16'b11111111_11001100;
   x93_i_tb = 16'b00000000_00010111;
   x94_r_tb = 16'b00000000_00111100;
   x94_i_tb = 16'b00000000_00011000;
   x95_r_tb = 16'b11111111_11000111;
   x95_i_tb = 16'b00000000_00010111; 
    x96_r_tb = 16'b11111111_11011011;
x96_i_tb =16'b11111111_11110000;
x97_r_tb = 16'b11111111_11011011;
x97_i_tb =16'b11111111_11110000;
x98_r_tb = 16'b11111111_11011011;
x98_i_tb =16'b11111111_11110000;
x99_r_tb = 16'b11111111_11011011;
x99_i_tb =16'b11111111_11110000;
x100_r_tb = 16'b11111111_11011011;
x100_i_tb =16'b11111111_11110000;
x101_r_tb = 16'b11111111_11011011;
x101_i_tb =16'b11111111_11110000;
x102_r_tb = 16'b11111111_11011011;
x102_i_tb =16'b11111111_11110000;
x103_r_tb = 16'b11111111_11011011;
x103_i_tb =16'b11111111_11110000;
x104_r_tb = 16'b11111111_11011011;
x104_i_tb =16'b11111111_11110000;
    x105_r_tb = 16'b11111111_11100010;
   x105_i_tb = 16'b00000000_00010100;
   x106_r_tb = 16'b00000000_00100010;
   x106_i_tb = 16'b00000000_00010100;
   x107_r_tb = 16'b11111111_11011011;
   x107_i_tb = 16'b11111111_11101011;
   x108_r_tb = 16'b00000000_00100110;
   x108_i_tb = 16'b11111111_11101011;
   x109_r_tb = 16'b11111111_11011000;
   x109_i_tb = 16'b00000000_00010011;
   x110_r_tb = 16'b00000000_00100111;
   x110_i_tb = 16'b00000000_00010001;
   x111_r_tb = 16'b00000000_00101000;
   x111_i_tb = 16'b00000000_00010001;
   x112_r_tb = 16'b11111111_11010100;
   x112_i_tb = 16'b11111111_11110000;
   x113_r_tb = 16'b00000000_00101110;
   x113_i_tb = 16'b11111111_11110010;
   x114_r_tb = 16'b11111111_11010001;
   x114_i_tb = 16'b00000000_00001100;
   x115_r_tb = 16'b00000000_00101011;
   x115_i_tb = 16'b00000000_00001100;
   x116_r_tb = 16'b00000000_00100111;
   x116_i_tb = 16'b00000000_00001010;
   x117_r_tb = 16'b11111111_11010100;
   x117_i_tb = 16'b00000000_00001010;
   x118_r_tb = 16'b11111111_11010010;
   x118_i_tb = 16'b11111111_11110010;
   x119_r_tb = 16'b00000000_00110000;
   x119_i_tb = 16'b11111111_11101101;
   x120_r_tb = 16'b11111111_11010010;
   x120_i_tb = 16'b00000000_00010100;
   x121_r_tb = 16'b00000000_00100111;
   x121_i_tb = 16'b11111111_11101011;
   x122_r_tb = 16'b00000000_00100010;
   x122_i_tb = 16'b00000000_00010001;
   x123_r_tb = 16'b00000000_00100111;
   x123_i_tb = 16'b00000000_00010100;
   x124_r_tb = 16'b00000000_00110000;
   x124_i_tb = 16'b11111111_11101100;
   x125_r_tb = 16'b11111111_11001100;
   x125_i_tb = 16'b00000000_00010111;
   x126_r_tb = 16'b00000000_00111100;
   x126_i_tb = 16'b00000000_00011000;
   x127_r_tb = 16'b11111111_11000111;
   x127_i_tb = 16'b00000000_00010111; 
 
   ready_inputs_tb = 1'b1 ;
    #(4*Clock_Period)
    ready_inputs_tb = 1'b0 ;


  end
endtask

   
endmodule

