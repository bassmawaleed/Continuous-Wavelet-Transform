module Reg_File #(

parameter NUMBER_OF_REGISTERS = 128 ,
parameter BITS = 16
)
( 
	input wire    [NUMBER_OF_REGISTERS - 1 : 0] WrEn , 
	input wire    clk ,
	input wire    rst , 

	input wire [BITS - 1 : 0] WrData_0,
	input wire [BITS - 1 : 0] WrData_1,
	input wire [BITS - 1 : 0] WrData_2,
	input wire [BITS - 1 : 0] WrData_3,
	input wire [BITS - 1 : 0] WrData_4,
	input wire [BITS - 1 : 0] WrData_5,
	input wire [BITS - 1 : 0] WrData_6,
	input wire [BITS - 1 : 0] WrData_7,
	input wire [BITS - 1 : 0] WrData_8,
	input wire [BITS - 1 : 0] WrData_9,
	input wire [BITS - 1 : 0] WrData_10,
	input wire [BITS - 1 : 0] WrData_11,
	input wire [BITS - 1 : 0] WrData_12,
	input wire [BITS - 1 : 0] WrData_13,
	input wire [BITS - 1 : 0] WrData_14,
	input wire [BITS - 1 : 0] WrData_15,
	input wire [BITS - 1 : 0] WrData_16,
	input wire [BITS - 1 : 0] WrData_17,
	input wire [BITS - 1 : 0] WrData_18,
	input wire [BITS - 1 : 0] WrData_19,
	input wire [BITS - 1 : 0] WrData_20,
	input wire [BITS - 1 : 0] WrData_21,
	input wire [BITS - 1 : 0] WrData_22,
	input wire [BITS - 1 : 0] WrData_23,
	input wire [BITS - 1 : 0] WrData_24,
	input wire [BITS - 1 : 0] WrData_25,
	input wire [BITS - 1 : 0] WrData_26,
	input wire [BITS - 1 : 0] WrData_27,
	input wire [BITS - 1 : 0] WrData_28,
	input wire [BITS - 1 : 0] WrData_29,
	input wire [BITS - 1 : 0] WrData_30,
	input wire [BITS - 1 : 0] WrData_31,
	input wire [BITS - 1 : 0] WrData_32,
	input wire [BITS - 1 : 0] WrData_33,
	input wire [BITS - 1 : 0] WrData_34,
	input wire [BITS - 1 : 0] WrData_35,
	input wire [BITS - 1 : 0] WrData_36,
	input wire [BITS - 1 : 0] WrData_37,
	input wire [BITS - 1 : 0] WrData_38,
	input wire [BITS - 1 : 0] WrData_39,
	input wire [BITS - 1 : 0] WrData_40,
	input wire [BITS - 1 : 0] WrData_41,
	input wire [BITS - 1 : 0] WrData_42,
	input wire [BITS - 1 : 0] WrData_43,
	input wire [BITS - 1 : 0] WrData_44,
	input wire [BITS - 1 : 0] WrData_45,
	input wire [BITS - 1 : 0] WrData_46,
	input wire [BITS - 1 : 0] WrData_47,
	input wire [BITS - 1 : 0] WrData_48,
	input wire [BITS - 1 : 0] WrData_49,
	input wire [BITS - 1 : 0] WrData_50,
	input wire [BITS - 1 : 0] WrData_51,
	input wire [BITS - 1 : 0] WrData_52,
	input wire [BITS - 1 : 0] WrData_53,
	input wire [BITS - 1 : 0] WrData_54,
	input wire [BITS - 1 : 0] WrData_55,
	input wire [BITS - 1 : 0] WrData_56,
	input wire [BITS - 1 : 0] WrData_57,
	input wire [BITS - 1 : 0] WrData_58,
	input wire [BITS - 1 : 0] WrData_59,
	input wire [BITS - 1 : 0] WrData_60,
	input wire [BITS - 1 : 0] WrData_61,
	input wire [BITS - 1 : 0] WrData_62,
	input wire [BITS - 1 : 0] WrData_63,
	input wire [BITS - 1 : 0] WrData_64,
	input wire [BITS - 1 : 0] WrData_65,
	input wire [BITS - 1 : 0] WrData_66,
	input wire [BITS - 1 : 0] WrData_67,
	input wire [BITS - 1 : 0] WrData_68,
	input wire [BITS - 1 : 0] WrData_69,
	input wire [BITS - 1 : 0] WrData_70,
	input wire [BITS - 1 : 0] WrData_71,
	input wire [BITS - 1 : 0] WrData_72,
	input wire [BITS - 1 : 0] WrData_73,
	input wire [BITS - 1 : 0] WrData_74,
	input wire [BITS - 1 : 0] WrData_75,
	input wire [BITS - 1 : 0] WrData_76,
	input wire [BITS - 1 : 0] WrData_77,
	input wire [BITS - 1 : 0] WrData_78,
	input wire [BITS - 1 : 0] WrData_79,
	input wire [BITS - 1 : 0] WrData_80,
	input wire [BITS - 1 : 0] WrData_81,
	input wire [BITS - 1 : 0] WrData_82,
	input wire [BITS - 1 : 0] WrData_83,
	input wire [BITS - 1 : 0] WrData_84,
	input wire [BITS - 1 : 0] WrData_85,
	input wire [BITS - 1 : 0] WrData_86,
	input wire [BITS - 1 : 0] WrData_87,
	input wire [BITS - 1 : 0] WrData_88,
	input wire [BITS - 1 : 0] WrData_89,
	input wire [BITS - 1 : 0] WrData_90,
	input wire [BITS - 1 : 0] WrData_91,
	input wire [BITS - 1 : 0] WrData_92,
	input wire [BITS - 1 : 0] WrData_93,
	input wire [BITS - 1 : 0] WrData_94,
	input wire [BITS - 1 : 0] WrData_95,
	input wire [BITS - 1 : 0] WrData_96,
	input wire [BITS - 1 : 0] WrData_97,
	input wire [BITS - 1 : 0] WrData_98,
	input wire [BITS - 1 : 0] WrData_99,
	input wire [BITS - 1 : 0] WrData_100,
	input wire [BITS - 1 : 0] WrData_101,
	input wire [BITS - 1 : 0] WrData_102,
	input wire [BITS - 1 : 0] WrData_103,
	input wire [BITS - 1 : 0] WrData_104,
	input wire [BITS - 1 : 0] WrData_105,
	input wire [BITS - 1 : 0] WrData_106,
	input wire [BITS - 1 : 0] WrData_107,
	input wire [BITS - 1 : 0] WrData_108,
	input wire [BITS - 1 : 0] WrData_109,
	input wire [BITS - 1 : 0] WrData_110,
	input wire [BITS - 1 : 0] WrData_111,
	input wire [BITS - 1 : 0] WrData_112,
	input wire [BITS - 1 : 0] WrData_113,
	input wire [BITS - 1 : 0] WrData_114,
	input wire [BITS - 1 : 0] WrData_115,
	input wire [BITS - 1 : 0] WrData_116,
	input wire [BITS - 1 : 0] WrData_117,
	input wire [BITS - 1 : 0] WrData_118,
	input wire [BITS - 1 : 0] WrData_119,
	input wire [BITS - 1 : 0] WrData_120,
	input wire [BITS - 1 : 0] WrData_121,
	input wire [BITS - 1 : 0] WrData_122,
	input wire [BITS - 1 : 0] WrData_123,
	input wire [BITS - 1 : 0] WrData_124,
	input wire [BITS - 1 : 0] WrData_125,
	input wire [BITS - 1 : 0] WrData_126,
	input wire [BITS - 1 : 0] WrData_127,



	output reg [BITS - 1 : 0] RdData_0,
	output reg [BITS - 1 : 0] RdData_1,
	output reg [BITS - 1 : 0] RdData_2,
	output reg [BITS - 1 : 0] RdData_3,
	output reg [BITS - 1 : 0] RdData_4,
	output reg [BITS - 1 : 0] RdData_5,
	output reg [BITS - 1 : 0] RdData_6,
	output reg [BITS - 1 : 0] RdData_7,
	output reg [BITS - 1 : 0] RdData_8,
	output reg [BITS - 1 : 0] RdData_9,
	output reg [BITS - 1 : 0] RdData_10,
	output reg [BITS - 1 : 0] RdData_11,
	output reg [BITS - 1 : 0] RdData_12,
	output reg [BITS - 1 : 0] RdData_13,
	output reg [BITS - 1 : 0] RdData_14,
	output reg [BITS - 1 : 0] RdData_15,
	output reg [BITS - 1 : 0] RdData_16,
	output reg [BITS - 1 : 0] RdData_17,
	output reg [BITS - 1 : 0] RdData_18,
	output reg [BITS - 1 : 0] RdData_19,
	output reg [BITS - 1 : 0] RdData_20,
	output reg [BITS - 1 : 0] RdData_21,
	output reg [BITS - 1 : 0] RdData_22,
	output reg [BITS - 1 : 0] RdData_23,
	output reg [BITS - 1 : 0] RdData_24,
	output reg [BITS - 1 : 0] RdData_25,
	output reg [BITS - 1 : 0] RdData_26,
	output reg [BITS - 1 : 0] RdData_27,
	output reg [BITS - 1 : 0] RdData_28,
	output reg [BITS - 1 : 0] RdData_29,
	output reg [BITS - 1 : 0] RdData_30,
	output reg [BITS - 1 : 0] RdData_31,
	output reg [BITS - 1 : 0] RdData_32,
	output reg [BITS - 1 : 0] RdData_33,
	output reg [BITS - 1 : 0] RdData_34,
	output reg [BITS - 1 : 0] RdData_35,
	output reg [BITS - 1 : 0] RdData_36,
	output reg [BITS - 1 : 0] RdData_37,
	output reg [BITS - 1 : 0] RdData_38,
	output reg [BITS - 1 : 0] RdData_39,
	output reg [BITS - 1 : 0] RdData_40,
	output reg [BITS - 1 : 0] RdData_41,
	output reg [BITS - 1 : 0] RdData_42,
	output reg [BITS - 1 : 0] RdData_43,
	output reg [BITS - 1 : 0] RdData_44,
	output reg [BITS - 1 : 0] RdData_45,
	output reg [BITS - 1 : 0] RdData_46,
	output reg [BITS - 1 : 0] RdData_47,
	output reg [BITS - 1 : 0] RdData_48,
	output reg [BITS - 1 : 0] RdData_49,
	output reg [BITS - 1 : 0] RdData_50,
	output reg [BITS - 1 : 0] RdData_51,
	output reg [BITS - 1 : 0] RdData_52,
	output reg [BITS - 1 : 0] RdData_53,
	output reg [BITS - 1 : 0] RdData_54,
	output reg [BITS - 1 : 0] RdData_55,
	output reg [BITS - 1 : 0] RdData_56,
	output reg [BITS - 1 : 0] RdData_57,
	output reg [BITS - 1 : 0] RdData_58,
	output reg [BITS - 1 : 0] RdData_59,
	output reg [BITS - 1 : 0] RdData_60,
	output reg [BITS - 1 : 0] RdData_61,
	output reg [BITS - 1 : 0] RdData_62,
	output reg [BITS - 1 : 0] RdData_63,
	output reg [BITS - 1 : 0] RdData_64,
	output reg [BITS - 1 : 0] RdData_65,
	output reg [BITS - 1 : 0] RdData_66,
	output reg [BITS - 1 : 0] RdData_67,
	output reg [BITS - 1 : 0] RdData_68,
	output reg [BITS - 1 : 0] RdData_69,
	output reg [BITS - 1 : 0] RdData_70,
	output reg [BITS - 1 : 0] RdData_71,
	output reg [BITS - 1 : 0] RdData_72,
	output reg [BITS - 1 : 0] RdData_73,
	output reg [BITS - 1 : 0] RdData_74,
	output reg [BITS - 1 : 0] RdData_75,
	output reg [BITS - 1 : 0] RdData_76,
	output reg [BITS - 1 : 0] RdData_77,
	output reg [BITS - 1 : 0] RdData_78,
	output reg [BITS - 1 : 0] RdData_79,
	output reg [BITS - 1 : 0] RdData_80,
	output reg [BITS - 1 : 0] RdData_81,
	output reg [BITS - 1 : 0] RdData_82,
	output reg [BITS - 1 : 0] RdData_83,
	output reg [BITS - 1 : 0] RdData_84,
	output reg [BITS - 1 : 0] RdData_85,
	output reg [BITS - 1 : 0] RdData_86,
	output reg [BITS - 1 : 0] RdData_87,
	output reg [BITS - 1 : 0] RdData_88,
	output reg [BITS - 1 : 0] RdData_89,
	output reg [BITS - 1 : 0] RdData_90,
	output reg [BITS - 1 : 0] RdData_91,
	output reg [BITS - 1 : 0] RdData_92,
	output reg [BITS - 1 : 0] RdData_93,
	output reg [BITS - 1 : 0] RdData_94,
	output reg [BITS - 1 : 0] RdData_95,
	output reg [BITS - 1 : 0] RdData_96,
	output reg [BITS - 1 : 0] RdData_97,
	output reg [BITS - 1 : 0] RdData_98,
	output reg [BITS - 1 : 0] RdData_99,
	output reg [BITS - 1 : 0] RdData_100,
	output reg [BITS - 1 : 0] RdData_101,
	output reg [BITS - 1 : 0] RdData_102,
	output reg [BITS - 1 : 0] RdData_103,
	output reg [BITS - 1 : 0] RdData_104,
	output reg [BITS - 1 : 0] RdData_105,
	output reg [BITS - 1 : 0] RdData_106,
	output reg [BITS - 1 : 0] RdData_107,
	output reg [BITS - 1 : 0] RdData_108,
	output reg [BITS - 1 : 0] RdData_109,
	output reg [BITS - 1 : 0] RdData_110,
	output reg [BITS - 1 : 0] RdData_111,
	output reg [BITS - 1 : 0] RdData_112,
	output reg [BITS - 1 : 0] RdData_113,
	output reg [BITS - 1 : 0] RdData_114,
	output reg [BITS - 1 : 0] RdData_115,
	output reg [BITS - 1 : 0] RdData_116,
	output reg [BITS - 1 : 0] RdData_117,
	output reg [BITS - 1 : 0] RdData_118,
	output reg [BITS - 1 : 0] RdData_119,
	output reg [BITS - 1 : 0] RdData_120,
	output reg [BITS - 1 : 0] RdData_121,
	output reg [BITS - 1 : 0] RdData_122,
	output reg [BITS - 1 : 0] RdData_123,
	output reg [BITS - 1 : 0] RdData_124,
	output reg [BITS - 1 : 0] RdData_125,
	output reg [BITS - 1 : 0] RdData_126,
	output reg [BITS - 1 : 0] RdData_127

  
  );
 
/* For Loop Counter */
integer i ;


always @ (posedge clk or negedge rst)
begin
  if ( !rst )
    begin
		RdData_0  <= 'b0;   RdData_1  <= 'b0;   RdData_2  <= 'b0;   RdData_3  <= 'b0;   RdData_4  <= 'b0;   RdData_5  <= 'b0;
		RdData_6  <= 'b0;   RdData_7  <= 'b0;   RdData_8  <= 'b0;   RdData_9  <= 'b0;   RdData_10 <= 'b0;   RdData_11 <= 'b0;
		RdData_12 <= 'b0;   RdData_13 <= 'b0;   RdData_14 <= 'b0;   RdData_15 <= 'b0;   RdData_16 <= 'b0;   RdData_17 <= 'b0;
		RdData_18 <= 'b0;   RdData_19 <= 'b0;   RdData_20 <= 'b0;   RdData_21 <= 'b0;   RdData_22 <= 'b0;   RdData_23 <= 'b0;
		RdData_24 <= 'b0;   RdData_25 <= 'b0;   RdData_26 <= 'b0;   RdData_27 <= 'b0;   RdData_28 <= 'b0;   RdData_29 <= 'b0;
		RdData_30 <= 'b0;   RdData_31 <= 'b0;   RdData_32 <= 'b0;   RdData_33 <= 'b0;   RdData_34 <= 'b0;   RdData_35 <= 'b0;
		RdData_36 <= 'b0;   RdData_37 <= 'b0;   RdData_38 <= 'b0;   RdData_39 <= 'b0;   RdData_40 <= 'b0;   RdData_41 <= 'b0;
		RdData_42 <= 'b0;   RdData_43 <= 'b0;   RdData_44 <= 'b0;   RdData_45 <= 'b0;   RdData_46 <= 'b0;   RdData_47 <= 'b0;
		RdData_48 <= 'b0;   RdData_49 <= 'b0;   RdData_50 <= 'b0;   RdData_51 <= 'b0;   RdData_52 <= 'b0;   RdData_53 <= 'b0;
		RdData_54 <= 'b0;   RdData_55 <= 'b0;

		RdData_56 <= 'b0;   RdData_57 <= 'b0;   RdData_58 <= 'b0;   RdData_59 <= 'b0;   RdData_60 <= 'b0;   RdData_61 <= 'b0;
		RdData_62 <= 'b0;   RdData_63 <= 'b0;   RdData_64 <= 'b0;   RdData_65 <= 'b0;   RdData_66 <= 'b0;   RdData_67 <= 'b0;
		RdData_68 <= 'b0;   RdData_69 <= 'b0;   RdData_70 <= 'b0;   RdData_71 <= 'b0;   RdData_72 <= 'b0;   RdData_73 <= 'b0;
		RdData_74 <= 'b0;   RdData_75 <= 'b0;   RdData_76 <= 'b0;   RdData_77 <= 'b0;   RdData_78 <= 'b0;   RdData_79 <= 'b0;
		RdData_80 <= 'b0;   RdData_81 <= 'b0;   RdData_82 <= 'b0;   RdData_83 <= 'b0;   RdData_84 <= 'b0;   RdData_85 <= 'b0;
		RdData_86 <= 'b0;   RdData_87 <= 'b0;   RdData_88 <= 'b0;   RdData_89 <= 'b0;   RdData_90 <= 'b0;   RdData_91 <= 'b0;
		RdData_92 <= 'b0;   RdData_93 <= 'b0;   RdData_94 <= 'b0;   RdData_95 <= 'b0;   RdData_96 <= 'b0;   RdData_97 <= 'b0;
		RdData_98 <= 'b0;   RdData_99 <= 'b0;   RdData_100 <= 'b0;  RdData_101 <= 'b0;  RdData_102 <= 'b0;  RdData_103 <= 'b0;
		RdData_104 <= 'b0;  RdData_105 <= 'b0;  RdData_106 <= 'b0;  RdData_107 <= 'b0;  RdData_108 <= 'b0;  RdData_109 <= 'b0;
		RdData_110 <= 'b0;  RdData_111 <= 'b0;

		RdData_112 <= 'b0;  RdData_113 <= 'b0;  RdData_114 <= 'b0;  RdData_115 <= 'b0;  RdData_116 <= 'b0;  RdData_117 <= 'b0;
		RdData_118 <= 'b0;  RdData_119 <= 'b0;  RdData_120 <= 'b0;  RdData_121 <= 'b0;  RdData_122 <= 'b0;  RdData_123 <= 'b0;
		RdData_124 <= 'b0;  RdData_125 <= 'b0;  RdData_126 <= 'b0;  RdData_127 <= 'b0; 
    end
  else
    begin
		if(WrEn[0] == 1)
		begin
			RdData_0 <= WrData_0 ;
		end
		
		if(WrEn[1] == 1)
		begin
			RdData_1 <= WrData_1 ;
		end
		
		if(WrEn[2] == 1)
		begin
			RdData_2 <= WrData_2 ;
		end
		
		if(WrEn[3] == 1)
		begin
			RdData_3 <= WrData_3 ;
		end
		
		if(WrEn[4] == 1)
		begin
			RdData_4 <= WrData_4 ;
		end
		
		if(WrEn[5] == 1)
		begin
			RdData_5 <= WrData_5 ;
		end
		
		if(WrEn[6] == 1)
		begin
			RdData_6 <= WrData_6 ;
		end
		
		if(WrEn[7] == 1)
		begin
			RdData_7 <= WrData_7 ;
		end
		
		if(WrEn[8] == 1)
		begin
			RdData_8 <= WrData_8 ;
		end
		
		if(WrEn[9] == 1)
		begin
			RdData_9 <= WrData_9 ;
		end
		
		if(WrEn[10] == 1)
		begin
			RdData_10 <= WrData_10 ;
		end
		
		if(WrEn[11] == 1)
		begin
			RdData_11 <= WrData_11 ;
		end
		
		if(WrEn[12] == 1)
		begin
			RdData_12 <= WrData_12 ;
		end
		
		if(WrEn[13] == 1)
		begin
			RdData_13 <= WrData_13 ;
		end
		
		if(WrEn[14] == 1)
		begin
			RdData_14 <= WrData_14 ;
		end
		
		if(WrEn[15] == 1)
		begin
			RdData_15 <= WrData_15 ;
		end
		
		if(WrEn[16] == 1)
		begin
			RdData_16 <= WrData_16 ;
		end
		
		if(WrEn[17] == 1)
		begin
			RdData_17 <= WrData_17 ;
		end
		
		if(WrEn[18] == 1)
		begin
			RdData_18 <= WrData_18 ;
		end
		
		if(WrEn[19] == 1)
		begin
			RdData_19 <= WrData_19 ;
		end
		
		if(WrEn[20] == 1)
		begin
			RdData_20 <= WrData_20 ;
		end
		
		if(WrEn[21] == 1)
		begin
			RdData_21 <= WrData_21 ;
		end
		
		if(WrEn[22] == 1)
		begin
			RdData_22 <= WrData_22 ;
		end
		
		if(WrEn[23] == 1)
		begin
			RdData_23 <= WrData_23 ;
		end
		
		if(WrEn[24] == 1)
		begin
			RdData_24 <= WrData_24 ;
		end
		
		if(WrEn[25] == 1)
		begin
			RdData_25 <= WrData_25 ;
		end
		
		if(WrEn[26] == 1)
		begin
			RdData_26 <= WrData_26 ;
		end
		
		if(WrEn[27] == 1)
		begin
			RdData_27 <= WrData_27 ;
		end
		
		if(WrEn[28] == 1)
		begin
			RdData_28 <= WrData_28 ;
		end
		
		if(WrEn[29] == 1)
		begin
			RdData_29 <= WrData_29 ;
		end
		
		if(WrEn[30] == 1)
		begin
			RdData_30 <= WrData_30 ;
		end
		
		if(WrEn[31] == 1)
		begin
			RdData_31 <= WrData_31 ;
		end
		
		if(WrEn[32] == 1)
		begin
			RdData_32 <= WrData_32 ;
		end
		
		if(WrEn[33] == 1)
		begin
			RdData_33 <= WrData_33 ;
		end
		
		if(WrEn[34] == 1)
		begin
			RdData_34 <= WrData_34 ;
		end
		
		if(WrEn[35] == 1)
		begin
			RdData_35 <= WrData_35 ;
		end
		
		if(WrEn[36] == 1)
		begin
			RdData_36 <= WrData_36 ;
		end
		
		if(WrEn[37] == 1)
		begin
			RdData_37 <= WrData_37 ;
		end
		
		if(WrEn[38] == 1)
		begin
			RdData_38 <= WrData_38 ;
		end
		
		if(WrEn[39] == 1)
		begin
			RdData_39 <= WrData_39 ;
		end
		
		if(WrEn[40] == 1)
		begin
			RdData_40 <= WrData_40 ;
		end
		
		if(WrEn[41] == 1)
		begin
			RdData_41 <= WrData_41 ;
		end
		
		if(WrEn[42] == 1)
		begin
			RdData_42 <= WrData_42 ;
		end
		
		if(WrEn[43] == 1)
		begin
			RdData_43 <= WrData_43 ;
		end
		
		if(WrEn[44] == 1)
		begin
			RdData_44 <= WrData_44 ;
		end
		
		if(WrEn[45] == 1)
		begin
			RdData_45 <= WrData_45 ;
		end
		
		if(WrEn[46] == 1)
		begin
			RdData_46 <= WrData_46 ;
		end
		
		if(WrEn[47] == 1)
		begin
			RdData_47 <= WrData_47 ;
		end
		
		if(WrEn[48] == 1)
		begin
			RdData_48 <= WrData_48 ;
		end
		
		if(WrEn[49] == 1)
		begin
			RdData_49 <= WrData_49 ;
		end
		
		if(WrEn[50] == 1)
		begin
			RdData_50 <= WrData_50 ;
		end
		
		if(WrEn[51] == 1)
		begin
			RdData_51 <= WrData_51 ;
		end
		
		if(WrEn[52] == 1)
		begin
			RdData_52 <= WrData_52 ;
		end
		
		if(WrEn[53] == 1)
		begin
			RdData_53 <= WrData_53 ;
		end
		
		if(WrEn[54] == 1)
		begin
			RdData_54 <= WrData_54 ;
		end
		
		if(WrEn[55] == 1)
		begin
			RdData_55 <= WrData_55 ;
		end
		
		if(WrEn[56] == 1)
		begin
			RdData_56 <= WrData_56 ;
		end
		
		if(WrEn[57] == 1)
		begin
			RdData_57 <= WrData_57 ;
		end
		
		if(WrEn[58] == 1)
		begin
			RdData_58 <= WrData_58 ;
		end
		
		if(WrEn[59] == 1)
		begin
			RdData_59 <= WrData_59 ;
		end
		
		if(WrEn[60] == 1)
		begin
			RdData_60 <= WrData_60 ;
		end
		
		if(WrEn[61] == 1)
		begin
			RdData_61 <= WrData_61 ;
		end
		
		if(WrEn[62] == 1)
		begin
			RdData_62 <= WrData_62 ;
		end
		
		if(WrEn[63] == 1)
		begin
			RdData_63 <= WrData_63 ;
		end
		
		if(WrEn[64] == 1)
		begin
			RdData_64 <= WrData_64 ;
		end
		
		if(WrEn[65] == 1)
		begin
			RdData_65 <= WrData_65 ;
		end
		
		if(WrEn[66] == 1)
		begin
			RdData_66 <= WrData_66 ;
		end
		
		if(WrEn[67] == 1)
		begin
			RdData_67 <= WrData_67 ;
		end
		
		if(WrEn[68] == 1)
		begin
			RdData_68 <= WrData_68 ;
		end
		
		if(WrEn[69] == 1)
		begin
			RdData_69 <= WrData_69 ;
		end
		
		if(WrEn[70] == 1)
		begin
			RdData_70 <= WrData_70 ;
		end
		
		if(WrEn[71] == 1)
		begin
			RdData_71 <= WrData_71 ;
		end
		
		if(WrEn[72] == 1)
		begin
			RdData_72 <= WrData_72 ;
		end
		
		if(WrEn[73] == 1)
		begin
			RdData_73 <= WrData_73 ;
		end
		
		if(WrEn[74] == 1)
		begin
			RdData_74 <= WrData_74 ;
		end
		
		if(WrEn[75] == 1)
		begin
			RdData_75 <= WrData_75 ;
		end
		
		if(WrEn[76] == 1)
		begin
			RdData_76 <= WrData_76 ;
		end
		
		if(WrEn[77] == 1)
		begin
			RdData_77 <= WrData_77 ;
		end
		
		if(WrEn[78] == 1)
		begin
			RdData_78 <= WrData_78 ;
		end
		
		if(WrEn[79] == 1)
		begin
			RdData_79 <= WrData_79 ;
		end
		
		if(WrEn[80] == 1)
		begin
			RdData_80 <= WrData_80 ;
		end
		
		if(WrEn[81] == 1)
		begin
			RdData_81 <= WrData_81 ;
		end
		
		if(WrEn[82] == 1)
		begin
			RdData_82 <= WrData_82 ;
		end
		
		if(WrEn[83] == 1)
		begin
			RdData_83 <= WrData_83 ;
		end
		
		if(WrEn[84] == 1)
		begin
			RdData_84 <= WrData_84 ;
		end
		
		if(WrEn[85] == 1)
		begin
			RdData_85 <= WrData_85 ;
		end
		
		if(WrEn[86] == 1)
		begin
			RdData_86 <= WrData_86 ;
		end
		
		if(WrEn[87] == 1)
		begin
			RdData_87 <= WrData_87 ;
		end
		
		if(WrEn[88] == 1)
		begin
			RdData_88 <= WrData_88 ;
		end
		
		if(WrEn[89] == 1)
		begin
			RdData_89 <= WrData_89 ;
		end
		
		if(WrEn[90] == 1)
		begin
			RdData_90 <= WrData_90 ;
		end
		
		if(WrEn[91] == 1)
		begin
			RdData_91 <= WrData_91 ;
		end
		
		if(WrEn[92] == 1)
		begin
			RdData_92 <= WrData_92 ;
		end
		
		if(WrEn[93] == 1)
		begin
			RdData_93 <= WrData_93 ;
		end
		
		if(WrEn[94] == 1)
		begin
			RdData_94 <= WrData_94 ;
		end
		
		if(WrEn[95] == 1)
		begin
			RdData_95 <= WrData_95 ;
		end
		
		if(WrEn[96] == 1)
		begin
			RdData_96 <= WrData_96 ;
		end
		
		if(WrEn[97] == 1)
		begin
			RdData_97 <= WrData_97 ;
		end
		
		if(WrEn[98] == 1)
		begin
			RdData_98 <= WrData_98 ;
		end
		
		if(WrEn[99] == 1)
		begin
			RdData_99 <= WrData_99 ;
		end
		
		if(WrEn[100] == 1)
		begin
			RdData_100 <= WrData_100 ;
		end
		
		if(WrEn[101] == 1)
		begin
			RdData_101 <= WrData_101 ;
		end
		
		if(WrEn[102] == 1)
		begin
			RdData_102 <= WrData_102 ;
		end
		
		if(WrEn[103] == 1)
		begin
			RdData_103 <= WrData_103 ;
		end
		
		if(WrEn[104] == 1)
		begin
			RdData_104 <= WrData_104 ;
		end
		
		if(WrEn[105] == 1)
		begin
			RdData_105 <= WrData_105 ;
		end
		
		if(WrEn[106] == 1)
		begin
			RdData_106 <= WrData_106 ;
		end
		
		if(WrEn[107] == 1)
		begin
			RdData_107 <= WrData_107 ;
		end
		
		if(WrEn[108] == 1)
		begin
			RdData_108 <= WrData_108 ;
		end
		
		if(WrEn[109] == 1)
		begin
			RdData_109 <= WrData_109 ;
		end
		
		if(WrEn[110] == 1)
		begin
			RdData_110 <= WrData_110 ;
		end
		
		if(WrEn[111] == 1)
		begin
			RdData_111 <= WrData_111 ;
		end
		
		if(WrEn[112] == 1)
		begin
			RdData_112 <= WrData_112 ;
		end
		
		if(WrEn[113] == 1)
		begin
			RdData_113 <= WrData_113 ;
		end
		
		if(WrEn[114] == 1)
		begin
			RdData_114 <= WrData_114 ;
		end
		
		if(WrEn[15] == 1)
		begin
			RdData_115 <= WrData_115 ;
		end
		
		if(WrEn[116] == 1)
		begin
			RdData_116 <= WrData_116 ;
		end
		
		if(WrEn[117] == 1)
		begin
			RdData_117 <= WrData_117 ;
		end
		
		if(WrEn[118] == 1)
		begin
			RdData_118 <= WrData_118 ;
		end
		
		if(WrEn[119] == 1)
		begin
			RdData_119 <= WrData_119 ;
		end
		
		if(WrEn[120] == 1)
		begin
			RdData_120 <= WrData_120 ;
		end
		
		if(WrEn[121] == 1)
		begin
			RdData_121 <= WrData_121 ;
		end
		
		if(WrEn[122] == 1)
		begin
			RdData_122 <= WrData_122 ;
		end
		
		if(WrEn[123] == 1)
		begin
			RdData_123 <= WrData_123 ;
		end
		
		if(WrEn[124] == 1)
		begin
			RdData_124 <= WrData_124 ;
		end
		
		if(WrEn[125] == 1)
		begin
			RdData_125 <= WrData_125 ;
		end
		
		if(WrEn[126] == 1)
		begin
			RdData_126 <= WrData_126 ;
		end
		
		if(WrEn[127] == 1)
		begin
			RdData_127 <= WrData_127 ;
		end
	end
end

endmodule
